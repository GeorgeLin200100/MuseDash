module ROM (
    input [11:0] addr,
    output reg [1:0] noteup,
    output reg [1:0] notedown
);

reg [3:0] ROM [0:4095];

initial begin
	ROM[0] = 4'b0000;
	ROM[1] = 4'b0000;
	ROM[2] = 4'b0000;
	ROM[3] = 4'b0000;
	ROM[4] = 4'b0000;
	ROM[5] = 4'b0000;
	ROM[6] = 4'b0000;
	ROM[7] = 4'b0000;
	ROM[8] = 4'b0000;
	ROM[9] = 4'b0000;
	ROM[10] = 4'b0000;
	ROM[11] = 4'b0000;
	ROM[12] = 4'b0000;
	ROM[13] = 4'b0000;
	ROM[14] = 4'b0000;
	ROM[15] = 4'b0000;
	ROM[16] = 4'b0000;
	ROM[17] = 4'b0000;
	ROM[18] = 4'b0000;
	ROM[19] = 4'b0000;
	ROM[20] = 4'b0000;
	ROM[21] = 4'b0000;
	ROM[22] = 4'b0000;
	ROM[23] = 4'b0000;
	ROM[24] = 4'b0000;
	ROM[25] = 4'b0000;
	ROM[26] = 4'b0000;
	ROM[27] = 4'b0000;
	ROM[28] = 4'b0000;
	ROM[29] = 4'b0000;
	ROM[30] = 4'b0000;
	ROM[31] = 4'b0000;
	ROM[32] = 4'b0000;
	ROM[33] = 4'b0000;
	ROM[34] = 4'b0000;
	ROM[35] = 4'b0000;
	ROM[36] = 4'b0000;
	ROM[37] = 4'b0000;
	ROM[38] = 4'b0000;
	ROM[39] = 4'b0000;
	ROM[40] = 4'b0000;
	ROM[41] = 4'b0000;
	ROM[42] = 4'b0000;
	ROM[43] = 4'b0000;
	ROM[44] = 4'b0000;
	ROM[45] = 4'b0000;
	ROM[46] = 4'b0000;
	ROM[47] = 4'b0000;
	ROM[48] = 4'b0000;
	ROM[49] = 4'b0000;
	ROM[50] = 4'b0000;
	ROM[51] = 4'b0000;
	ROM[52] = 4'b0000;
	ROM[53] = 4'b0000;
	ROM[54] = 4'b0000;
	ROM[55] = 4'b0000;
	ROM[56] = 4'b0000;
	ROM[57] = 4'b0000;
	ROM[58] = 4'b0000;
	ROM[59] = 4'b0000;
	ROM[60] = 4'b0000;
	ROM[61] = 4'b0000;
	ROM[62] = 4'b0000;
	ROM[63] = 4'b0000;
	ROM[64] = 4'b0000;
	ROM[65] = 4'b0001;
	ROM[66] = 4'b0000;
	ROM[67] = 4'b0000;
	ROM[68] = 4'b0000;
	ROM[69] = 4'b0000;
	ROM[70] = 4'b0000;
	ROM[71] = 4'b0000;
	ROM[72] = 4'b0000;
	ROM[73] = 4'b0001;
	ROM[74] = 4'b0000;
	ROM[75] = 4'b0000;
	ROM[76] = 4'b0000;
	ROM[77] = 4'b0000;
	ROM[78] = 4'b0000;
	ROM[79] = 4'b0000;
	ROM[80] = 4'b0000;
	ROM[81] = 4'b0001;
	ROM[82] = 4'b0000;
	ROM[83] = 4'b0000;
	ROM[84] = 4'b0000;
	ROM[85] = 4'b0000;
	ROM[86] = 4'b0000;
	ROM[87] = 4'b0000;
	ROM[88] = 4'b0000;
	ROM[89] = 4'b0001;
	ROM[90] = 4'b0000;
	ROM[91] = 4'b0000;
	ROM[92] = 4'b0000;
	ROM[93] = 4'b0000;
	ROM[94] = 4'b0000;
	ROM[95] = 4'b0000;
	ROM[96] = 4'b0000;
	ROM[97] = 4'b0100;
	ROM[98] = 4'b0000;
	ROM[99] = 4'b0000;
	ROM[100] = 4'b0000;
	ROM[101] = 4'b0000;
	ROM[102] = 4'b0000;
	ROM[103] = 4'b0000;
	ROM[104] = 4'b0000;
	ROM[105] = 4'b0100;
	ROM[106] = 4'b0000;
	ROM[107] = 4'b0000;
	ROM[108] = 4'b0000;
	ROM[109] = 4'b0000;
	ROM[110] = 4'b0000;
	ROM[111] = 4'b0000;
	ROM[112] = 4'b0000;
	ROM[113] = 4'b0100;
	ROM[114] = 4'b0000;
	ROM[115] = 4'b0000;
	ROM[116] = 4'b0000;
	ROM[117] = 4'b0000;
	ROM[118] = 4'b0000;
	ROM[119] = 4'b0000;
	ROM[120] = 4'b0000;
	ROM[121] = 4'b0100;
	ROM[122] = 4'b0000;
	ROM[123] = 4'b0000;
	ROM[124] = 4'b0000;
	ROM[125] = 4'b0000;
	ROM[126] = 4'b0000;
	ROM[127] = 4'b0000;
	ROM[128] = 4'b0000;
	ROM[129] = 4'b0001;
	ROM[130] = 4'b0000;
	ROM[131] = 4'b0000;
	ROM[132] = 4'b0000;
	ROM[133] = 4'b0000;
	ROM[134] = 4'b0000;
	ROM[135] = 4'b0000;
	ROM[136] = 4'b0000;
	ROM[137] = 4'b0001;
	ROM[138] = 4'b0000;
	ROM[139] = 4'b0000;
	ROM[140] = 4'b0000;
	ROM[141] = 4'b0000;
	ROM[142] = 4'b0000;
	ROM[143] = 4'b0000;
	ROM[144] = 4'b0000;
	ROM[145] = 4'b0001;
	ROM[146] = 4'b0000;
	ROM[147] = 4'b0000;
	ROM[148] = 4'b0000;
	ROM[149] = 4'b0000;
	ROM[150] = 4'b0000;
	ROM[151] = 4'b0000;
	ROM[152] = 4'b0000;
	ROM[153] = 4'b0001;
	ROM[154] = 4'b0000;
	ROM[155] = 4'b0000;
	ROM[156] = 4'b0000;
	ROM[157] = 4'b0000;
	ROM[158] = 4'b0000;
	ROM[159] = 4'b0000;
	ROM[160] = 4'b0000;
	ROM[161] = 4'b0100;
	ROM[162] = 4'b0000;
	ROM[163] = 4'b0000;
	ROM[164] = 4'b0000;
	ROM[165] = 4'b0000;
	ROM[166] = 4'b0000;
	ROM[167] = 4'b0000;
	ROM[168] = 4'b0000;
	ROM[169] = 4'b0100;
	ROM[170] = 4'b0000;
	ROM[171] = 4'b0000;
	ROM[172] = 4'b0000;
	ROM[173] = 4'b0000;
	ROM[174] = 4'b0000;
	ROM[175] = 4'b0000;
	ROM[176] = 4'b0000;
	ROM[177] = 4'b0100;
	ROM[178] = 4'b0000;
	ROM[179] = 4'b0000;
	ROM[180] = 4'b0000;
	ROM[181] = 4'b0100;
	ROM[182] = 4'b0000;
	ROM[183] = 4'b0000;
	ROM[184] = 4'b0000;
	ROM[185] = 4'b0100;
	ROM[186] = 4'b0000;
	ROM[187] = 4'b0100;
	ROM[188] = 4'b0000;
	ROM[189] = 4'b0100;
	ROM[190] = 4'b0000;
	ROM[191] = 4'b0000;
	ROM[192] = 4'b0000;
	ROM[193] = 4'b0001;
	ROM[194] = 4'b0000;
	ROM[195] = 4'b0001;
	ROM[196] = 4'b0000;
	ROM[197] = 4'b0001;
	ROM[198] = 4'b0000;
	ROM[199] = 4'b0001;
	ROM[200] = 4'b0000;
	ROM[201] = 4'b0100;
	ROM[202] = 4'b0000;
	ROM[203] = 4'b0100;
	ROM[204] = 4'b0000;
	ROM[205] = 4'b0100;
	ROM[206] = 4'b0000;
	ROM[207] = 4'b0100;
	ROM[208] = 4'b0000;
	ROM[209] = 4'b0001;
	ROM[210] = 4'b0000;
	ROM[211] = 4'b0000;
	ROM[212] = 4'b0001;
	ROM[213] = 4'b0000;
	ROM[214] = 4'b0000;
	ROM[215] = 4'b0001;
	ROM[216] = 4'b0000;
	ROM[217] = 4'b0001;
	ROM[218] = 4'b0000;
	ROM[219] = 4'b0000;
	ROM[220] = 4'b0000;
	ROM[221] = 4'b0100;
	ROM[222] = 4'b0000;
	ROM[223] = 4'b0000;
	ROM[224] = 4'b0000;
	ROM[225] = 4'b0001;
	ROM[226] = 4'b0000;
	ROM[227] = 4'b0000;
	ROM[228] = 4'b0000;
	ROM[229] = 4'b0100;
	ROM[230] = 4'b0000;
	ROM[231] = 4'b0000;
	ROM[232] = 4'b0000;
	ROM[233] = 4'b0001;
	ROM[234] = 4'b0000;
	ROM[235] = 4'b0000;
	ROM[236] = 4'b0000;
	ROM[237] = 4'b0100;
	ROM[238] = 4'b0000;
	ROM[239] = 4'b0000;
	ROM[240] = 4'b0000;
	ROM[241] = 4'b1000;
	ROM[242] = 4'b1100;
	ROM[243] = 4'b1100;
	ROM[244] = 4'b1100;
	ROM[245] = 4'b1100;
	ROM[246] = 4'b1100;
	ROM[247] = 4'b1100;
	ROM[248] = 4'b1100;
	ROM[249] = 4'b1100;
	ROM[250] = 4'b1100;
	ROM[251] = 4'b1100;
	ROM[252] = 4'b1100;
	ROM[253] = 4'b1100;
	ROM[254] = 4'b1100;
	ROM[255] = 4'b1100;
	ROM[256] = 4'b1100;
	ROM[257] = 4'b1110;
	ROM[258] = 4'b0011;
	ROM[259] = 4'b0011;
	ROM[260] = 4'b0011;
	ROM[261] = 4'b0111;
	ROM[262] = 4'b0000;
	ROM[263] = 4'b0100;
	ROM[264] = 4'b0000;
	ROM[265] = 4'b0001;
	ROM[266] = 4'b0000;
	ROM[267] = 4'b0001;
	ROM[268] = 4'b0000;
	ROM[269] = 4'b0100;
	ROM[270] = 4'b0000;
	ROM[271] = 4'b0100;
	ROM[272] = 4'b0000;
	ROM[273] = 4'b0001;
	ROM[274] = 4'b0000;
	ROM[275] = 4'b0001;
	ROM[276] = 4'b0000;
	ROM[277] = 4'b0100;
	ROM[278] = 4'b0000;
	ROM[279] = 4'b0100;
	ROM[280] = 4'b0000;
	ROM[281] = 4'b0001;
	ROM[282] = 4'b0000;
	ROM[283] = 4'b0010;
	ROM[284] = 4'b0011;
	ROM[285] = 4'b0011;
	ROM[286] = 4'b0011;
	ROM[287] = 4'b0111;
	ROM[288] = 4'b0000;
	ROM[289] = 4'b0100;
	ROM[290] = 4'b0000;
	ROM[291] = 4'b0001;
	ROM[292] = 4'b0000;
	ROM[293] = 4'b0010;
	ROM[294] = 4'b0011;
	ROM[295] = 4'b0011;
	ROM[296] = 4'b0011;
	ROM[297] = 4'b0111;
	ROM[298] = 4'b0000;
	ROM[299] = 4'b0100;
	ROM[300] = 4'b0000;
	ROM[301] = 4'b0001;
	ROM[302] = 4'b0000;
	ROM[303] = 4'b0001;
	ROM[304] = 4'b0000;
	ROM[305] = 4'b1000;
	ROM[306] = 4'b1100;
	ROM[307] = 4'b1100;
	ROM[308] = 4'b1100;
	ROM[309] = 4'b1100;
	ROM[310] = 4'b1100;
	ROM[311] = 4'b1100;
	ROM[312] = 4'b1100;
	ROM[313] = 4'b1110;
	ROM[314] = 4'b0011;
	ROM[315] = 4'b0011;
	ROM[316] = 4'b0011;
	ROM[317] = 4'b0011;
	ROM[318] = 4'b0011;
	ROM[319] = 4'b0011;
	ROM[320] = 4'b0011;
	ROM[321] = 4'b0111;
	ROM[322] = 4'b0000;
	ROM[323] = 4'b0000;
	ROM[324] = 4'b0000;
	ROM[325] = 4'b0000;
	ROM[326] = 4'b0000;
	ROM[327] = 4'b0000;
	ROM[328] = 4'b0000;
	ROM[329] = 4'b0000;
	ROM[330] = 4'b0000;
	ROM[331] = 4'b0000;
	ROM[332] = 4'b0000;
	ROM[333] = 4'b0000;
	ROM[334] = 4'b0000;
	ROM[335] = 4'b0000;
	ROM[336] = 4'b0000;
	ROM[337] = 4'b0001;
	ROM[338] = 4'b0000;
	ROM[339] = 4'b0000;
	ROM[340] = 4'b0000;
	ROM[341] = 4'b0001;
	ROM[342] = 4'b0000;
	ROM[343] = 4'b0001;
	ROM[344] = 4'b0000;
	ROM[345] = 4'b0001;
	ROM[346] = 4'b0000;
	ROM[347] = 4'b0000;
	ROM[348] = 4'b0000;
	ROM[349] = 4'b0100;
	ROM[350] = 4'b0000;
	ROM[351] = 4'b0000;
	ROM[352] = 4'b0000;
	ROM[353] = 4'b0001;
	ROM[354] = 4'b0000;
	ROM[355] = 4'b0000;
	ROM[356] = 4'b0000;
	ROM[357] = 4'b0101;
	ROM[358] = 4'b0000;
	ROM[359] = 4'b0000;
	ROM[360] = 4'b0000;
	ROM[361] = 4'b0001;
	ROM[362] = 4'b0000;
	ROM[363] = 4'b0000;
	ROM[364] = 4'b0000;
	ROM[365] = 4'b0101;
	ROM[366] = 4'b0000;
	ROM[367] = 4'b0000;
	ROM[368] = 4'b0000;
	ROM[369] = 4'b0100;
	ROM[370] = 4'b0000;
	ROM[371] = 4'b0000;
	ROM[372] = 4'b0000;
	ROM[373] = 4'b0101;
	ROM[374] = 4'b0000;
	ROM[375] = 4'b0000;
	ROM[376] = 4'b0000;
	ROM[377] = 4'b0100;
	ROM[378] = 4'b0000;
	ROM[379] = 4'b0000;
	ROM[380] = 4'b0000;
	ROM[381] = 4'b0101;
	ROM[382] = 4'b0000;
	ROM[383] = 4'b0000;
	ROM[384] = 4'b0000;
	ROM[385] = 4'b0001;
	ROM[386] = 4'b0000;
	ROM[387] = 4'b0000;
	ROM[388] = 4'b0000;
	ROM[389] = 4'b0101;
	ROM[390] = 4'b0000;
	ROM[391] = 4'b0000;
	ROM[392] = 4'b0000;
	ROM[393] = 4'b0001;
	ROM[394] = 4'b0000;
	ROM[395] = 4'b0000;
	ROM[396] = 4'b0000;
	ROM[397] = 4'b0101;
	ROM[398] = 4'b0000;
	ROM[399] = 4'b0000;
	ROM[400] = 4'b0000;
	ROM[401] = 4'b0100;
	ROM[402] = 4'b0000;
	ROM[403] = 4'b0000;
	ROM[404] = 4'b0000;
	ROM[405] = 4'b0101;
	ROM[406] = 4'b0000;
	ROM[407] = 4'b0000;
	ROM[408] = 4'b0000;
	ROM[409] = 4'b0100;
	ROM[410] = 4'b0000;
	ROM[411] = 4'b0000;
	ROM[412] = 4'b0000;
	ROM[413] = 4'b0101;
	ROM[414] = 4'b0000;
	ROM[415] = 4'b0000;
	ROM[416] = 4'b0000;
	ROM[417] = 4'b0001;
	ROM[418] = 4'b0000;
	ROM[419] = 4'b0001;
	ROM[420] = 4'b0000;
	ROM[421] = 4'b0100;
	ROM[422] = 4'b0000;
	ROM[423] = 4'b0100;
	ROM[424] = 4'b0000;
	ROM[425] = 4'b0001;
	ROM[426] = 4'b0000;
	ROM[427] = 4'b0001;
	ROM[428] = 4'b0000;
	ROM[429] = 4'b0100;
	ROM[430] = 4'b0000;
	ROM[431] = 4'b0100;
	ROM[432] = 4'b0000;
	ROM[433] = 4'b0001;
	ROM[434] = 4'b0000;
	ROM[435] = 4'b0000;
	ROM[436] = 4'b0001;
	ROM[437] = 4'b0000;
	ROM[438] = 4'b0000;
	ROM[439] = 4'b0001;
	ROM[440] = 4'b0000;
	ROM[441] = 4'b0001;
	ROM[442] = 4'b0000;
	ROM[443] = 4'b0000;
	ROM[444] = 4'b0000;
	ROM[445] = 4'b0100;
	ROM[446] = 4'b0000;
	ROM[447] = 4'b0000;
	ROM[448] = 4'b0000;
	ROM[449] = 4'b0001;
	ROM[450] = 4'b0000;
	ROM[451] = 4'b0001;
	ROM[452] = 4'b0000;
	ROM[453] = 4'b0100;
	ROM[454] = 4'b0000;
	ROM[455] = 4'b0100;
	ROM[456] = 4'b0000;
	ROM[457] = 4'b0001;
	ROM[458] = 4'b0000;
	ROM[459] = 4'b0001;
	ROM[460] = 4'b0000;
	ROM[461] = 4'b0100;
	ROM[462] = 4'b0000;
	ROM[463] = 4'b0100;
	ROM[464] = 4'b0000;
	ROM[465] = 4'b0001;
	ROM[466] = 4'b0000;
	ROM[467] = 4'b0000;
	ROM[468] = 4'b0000;
	ROM[469] = 4'b0001;
	ROM[470] = 4'b0000;
	ROM[471] = 4'b0000;
	ROM[472] = 4'b0000;
	ROM[473] = 4'b0001;
	ROM[474] = 4'b0000;
	ROM[475] = 4'b0000;
	ROM[476] = 4'b0000;
	ROM[477] = 4'b0100;
	ROM[478] = 4'b0000;
	ROM[479] = 4'b0000;
	ROM[480] = 4'b0000;
	ROM[481] = 4'b0001;
	ROM[482] = 4'b0000;
	ROM[483] = 4'b0001;
	ROM[484] = 4'b0000;
	ROM[485] = 4'b0000;
	ROM[486] = 4'b0000;
	ROM[487] = 4'b0100;
	ROM[488] = 4'b0000;
	ROM[489] = 4'b0100;
	ROM[490] = 4'b0000;
	ROM[491] = 4'b0000;
	ROM[492] = 4'b0000;
	ROM[493] = 4'b0001;
	ROM[494] = 4'b0000;
	ROM[495] = 4'b0001;
	ROM[496] = 4'b0000;
	ROM[497] = 4'b0000;
	ROM[498] = 4'b0000;
	ROM[499] = 4'b0100;
	ROM[500] = 4'b0000;
	ROM[501] = 4'b0100;
	ROM[502] = 4'b0000;
	ROM[503] = 4'b0000;
	ROM[504] = 4'b0000;
	ROM[505] = 4'b0001;
	ROM[506] = 4'b0000;
	ROM[507] = 4'b0000;
	ROM[508] = 4'b0000;
	ROM[509] = 4'b0100;
	ROM[510] = 4'b0000;
	ROM[511] = 4'b0000;
	ROM[512] = 4'b0000;
	ROM[513] = 4'b0001;
	ROM[514] = 4'b0000;
	ROM[515] = 4'b0000;
	ROM[516] = 4'b0000;
	ROM[517] = 4'b0100;
	ROM[518] = 4'b0000;
	ROM[519] = 4'b0000;
	ROM[520] = 4'b0000;
	ROM[521] = 4'b0001;
	ROM[522] = 4'b0000;
	ROM[523] = 4'b0001;
	ROM[524] = 4'b0000;
	ROM[525] = 4'b0000;
	ROM[526] = 4'b0000;
	ROM[527] = 4'b0100;
	ROM[528] = 4'b0000;
	ROM[529] = 4'b0001;
	ROM[530] = 4'b0000;
	ROM[531] = 4'b0000;
	ROM[532] = 4'b0000;
	ROM[533] = 4'b0001;
	ROM[534] = 4'b0000;
	ROM[535] = 4'b0000;
	ROM[536] = 4'b0000;
	ROM[537] = 4'b0100;
	ROM[538] = 4'b0000;
	ROM[539] = 4'b0100;
	ROM[540] = 4'b0000;
	ROM[541] = 4'b0100;
	ROM[542] = 4'b0000;
	ROM[543] = 4'b0000;
	ROM[544] = 4'b0000;
	ROM[545] = 4'b0001;
	ROM[546] = 4'b0000;
	ROM[547] = 4'b0001;
	ROM[548] = 4'b0000;
	ROM[549] = 4'b0000;
	ROM[550] = 4'b0000;
	ROM[551] = 4'b0100;
	ROM[552] = 4'b0000;
	ROM[553] = 4'b0100;
	ROM[554] = 4'b0000;
	ROM[555] = 4'b0000;
	ROM[556] = 4'b0000;
	ROM[557] = 4'b0001;
	ROM[558] = 4'b0000;
	ROM[559] = 4'b0001;
	ROM[560] = 4'b0000;
	ROM[561] = 4'b0000;
	ROM[562] = 4'b0000;
	ROM[563] = 4'b0100;
	ROM[564] = 4'b0000;
	ROM[565] = 4'b0100;
	ROM[566] = 4'b0000;
	ROM[567] = 4'b0000;
	ROM[568] = 4'b0000;
	ROM[569] = 4'b0001;
	ROM[570] = 4'b0000;
	ROM[571] = 4'b0000;
	ROM[572] = 4'b0000;
	ROM[573] = 4'b0100;
	ROM[574] = 4'b0000;
	ROM[575] = 4'b0000;
	ROM[576] = 4'b0000;
	ROM[577] = 4'b0001;
	ROM[578] = 4'b0000;
	ROM[579] = 4'b0000;
	ROM[580] = 4'b0000;
	ROM[581] = 4'b0100;
	ROM[582] = 4'b0000;
	ROM[583] = 4'b0000;
	ROM[584] = 4'b0000;
	ROM[585] = 4'b0001;
	ROM[586] = 4'b0000;
	ROM[587] = 4'b0001;
	ROM[588] = 4'b0000;
	ROM[589] = 4'b0000;
	ROM[590] = 4'b0000;
	ROM[591] = 4'b0100;
	ROM[592] = 4'b0000;
	ROM[593] = 4'b0001;
	ROM[594] = 4'b0000;
	ROM[595] = 4'b0000;
	ROM[596] = 4'b0000;
	ROM[597] = 4'b0001;
	ROM[598] = 4'b0000;
	ROM[599] = 4'b0000;
	ROM[600] = 4'b0000;
	ROM[601] = 4'b0001;
	ROM[602] = 4'b0000;
	ROM[603] = 4'b0000;
	ROM[604] = 4'b0000;
	ROM[605] = 4'b0100;
	ROM[606] = 4'b0000;
	ROM[607] = 4'b0000;
	ROM[608] = 4'b0000;
	ROM[609] = 4'b0001;
	ROM[610] = 4'b0000;
	ROM[611] = 4'b0001;
	ROM[612] = 4'b0000;
	ROM[613] = 4'b0100;
	ROM[614] = 4'b0000;
	ROM[615] = 4'b0001;
	ROM[616] = 4'b0000;
	ROM[617] = 4'b0001;
	ROM[618] = 4'b0000;
	ROM[619] = 4'b0000;
	ROM[620] = 4'b0000;
	ROM[621] = 4'b0100;
	ROM[622] = 4'b0000;
	ROM[623] = 4'b0100;
	ROM[624] = 4'b0000;
	ROM[625] = 4'b0001;
	ROM[626] = 4'b0000;
	ROM[627] = 4'b0100;
	ROM[628] = 4'b0000;
	ROM[629] = 4'b0100;
	ROM[630] = 4'b0000;
	ROM[631] = 4'b0000;
	ROM[632] = 4'b0000;
	ROM[633] = 4'b0001;
	ROM[634] = 4'b0000;
	ROM[635] = 4'b0000;
	ROM[636] = 4'b0000;
	ROM[637] = 4'b0100;
	ROM[638] = 4'b0000;
	ROM[639] = 4'b0000;
	ROM[640] = 4'b0000;
	ROM[641] = 4'b0001;
	ROM[642] = 4'b0000;
	ROM[643] = 4'b0000;
	ROM[644] = 4'b0000;
	ROM[645] = 4'b0100;
	ROM[646] = 4'b0000;
	ROM[647] = 4'b0000;
	ROM[648] = 4'b0000;
	ROM[649] = 4'b0001;
	ROM[650] = 4'b0000;
	ROM[651] = 4'b0001;
	ROM[652] = 4'b0000;
	ROM[653] = 4'b0100;
	ROM[654] = 4'b0000;
	ROM[655] = 4'b0001;
	ROM[656] = 4'b0000;
	ROM[657] = 4'b0100;
	ROM[658] = 4'b0000;
	ROM[659] = 4'b0100;
	ROM[660] = 4'b0000;
	ROM[661] = 4'b0001;
	ROM[662] = 4'b0000;
	ROM[663] = 4'b0001;
	ROM[664] = 4'b0000;
	ROM[665] = 4'b0100;
	ROM[666] = 4'b0000;
	ROM[667] = 4'b0100;
	ROM[668] = 4'b0000;
	ROM[669] = 4'b0001;
	ROM[670] = 4'b0000;
	ROM[671] = 4'b0001;
	ROM[672] = 4'b0000;
	ROM[673] = 4'b0100;
	ROM[674] = 4'b0000;
	ROM[675] = 4'b0100;
	ROM[676] = 4'b0000;
	ROM[677] = 4'b0001;
	ROM[678] = 4'b0000;
	ROM[679] = 4'b0100;
	ROM[680] = 4'b0000;
	ROM[681] = 4'b0000;
	ROM[682] = 4'b0000;
	ROM[683] = 4'b0001;
	ROM[684] = 4'b0000;
	ROM[685] = 4'b0001;
	ROM[686] = 4'b0000;
	ROM[687] = 4'b0000;
	ROM[688] = 4'b0000;
	ROM[689] = 4'b0100;
	ROM[690] = 4'b0000;
	ROM[691] = 4'b0001;
	ROM[692] = 4'b0000;
	ROM[693] = 4'b0100;
	ROM[694] = 4'b0000;
	ROM[695] = 4'b0000;
	ROM[696] = 4'b0000;
	ROM[697] = 4'b0001;
	ROM[698] = 4'b0000;
	ROM[699] = 4'b0100;
	ROM[700] = 4'b0000;
	ROM[701] = 4'b0001;
	ROM[702] = 4'b0000;
	ROM[703] = 4'b0000;
	ROM[704] = 4'b0000;
	ROM[705] = 4'b0100;
	ROM[706] = 4'b0000;
	ROM[707] = 4'b0100;
	ROM[708] = 4'b0000;
	ROM[709] = 4'b0100;
	ROM[710] = 4'b0000;
	ROM[711] = 4'b0000;
	ROM[712] = 4'b0000;
	ROM[713] = 4'b0001;
	ROM[714] = 4'b0000;
	ROM[715] = 4'b0001;
	ROM[716] = 4'b0000;
	ROM[717] = 4'b0001;
	ROM[718] = 4'b0000;
	ROM[719] = 4'b0000;
	ROM[720] = 4'b0000;
	ROM[721] = 4'b0100;
	ROM[722] = 4'b0000;
	ROM[723] = 4'b0000;
	ROM[724] = 4'b0100;
	ROM[725] = 4'b0000;
	ROM[726] = 4'b0000;
	ROM[727] = 4'b0001;
	ROM[728] = 4'b0000;
	ROM[729] = 4'b0001;
	ROM[730] = 4'b0000;
	ROM[731] = 4'b0000;
	ROM[732] = 4'b0000;
	ROM[733] = 4'b0100;
	ROM[734] = 4'b0000;
	ROM[735] = 4'b0000;
	ROM[736] = 4'b0000;
	ROM[737] = 4'b0001;
	ROM[738] = 4'b0000;
	ROM[739] = 4'b0001;
	ROM[740] = 4'b0000;
	ROM[741] = 4'b0100;
	ROM[742] = 4'b0000;
	ROM[743] = 4'b0001;
	ROM[744] = 4'b0000;
	ROM[745] = 4'b0001;
	ROM[746] = 4'b0000;
	ROM[747] = 4'b0000;
	ROM[748] = 4'b0000;
	ROM[749] = 4'b0100;
	ROM[750] = 4'b0000;
	ROM[751] = 4'b0100;
	ROM[752] = 4'b0000;
	ROM[753] = 4'b0001;
	ROM[754] = 4'b0000;
	ROM[755] = 4'b0100;
	ROM[756] = 4'b0000;
	ROM[757] = 4'b0100;
	ROM[758] = 4'b0000;
	ROM[759] = 4'b0000;
	ROM[760] = 4'b0000;
	ROM[761] = 4'b0001;
	ROM[762] = 4'b0000;
	ROM[763] = 4'b0000;
	ROM[764] = 4'b0000;
	ROM[765] = 4'b0100;
	ROM[766] = 4'b0000;
	ROM[767] = 4'b0000;
	ROM[768] = 4'b0000;
	ROM[769] = 4'b0001;
	ROM[770] = 4'b0000;
	ROM[771] = 4'b0000;
	ROM[772] = 4'b0000;
	ROM[773] = 4'b0100;
	ROM[774] = 4'b0000;
	ROM[775] = 4'b0000;
	ROM[776] = 4'b0000;
	ROM[777] = 4'b0001;
	ROM[778] = 4'b0000;
	ROM[779] = 4'b0001;
	ROM[780] = 4'b0000;
	ROM[781] = 4'b0100;
	ROM[782] = 4'b0000;
	ROM[783] = 4'b0001;
	ROM[784] = 4'b0000;
	ROM[785] = 4'b0100;
	ROM[786] = 4'b0000;
	ROM[787] = 4'b0100;
	ROM[788] = 4'b0000;
	ROM[789] = 4'b0001;
	ROM[790] = 4'b0000;
	ROM[791] = 4'b0001;
	ROM[792] = 4'b0000;
	ROM[793] = 4'b0100;
	ROM[794] = 4'b0000;
	ROM[795] = 4'b0100;
	ROM[796] = 4'b0000;
	ROM[797] = 4'b0001;
	ROM[798] = 4'b0000;
	ROM[799] = 4'b0001;
	ROM[800] = 4'b0000;
	ROM[801] = 4'b0100;
	ROM[802] = 4'b0000;
	ROM[803] = 4'b0100;
	ROM[804] = 4'b0000;
	ROM[805] = 4'b0001;
	ROM[806] = 4'b0000;
	ROM[807] = 4'b0100;
	ROM[808] = 4'b0000;
	ROM[809] = 4'b0000;
	ROM[810] = 4'b0000;
	ROM[811] = 4'b0001;
	ROM[812] = 4'b0000;
	ROM[813] = 4'b0001;
	ROM[814] = 4'b0000;
	ROM[815] = 4'b0000;
	ROM[816] = 4'b0000;
	ROM[817] = 4'b0100;
	ROM[818] = 4'b0000;
	ROM[819] = 4'b0000;
	ROM[820] = 4'b0000;
	ROM[821] = 4'b0001;
	ROM[822] = 4'b0000;
	ROM[823] = 4'b0000;
	ROM[824] = 4'b0000;
	ROM[825] = 4'b0100;
	ROM[826] = 4'b0000;
	ROM[827] = 4'b0000;
	ROM[828] = 4'b0000;
	ROM[829] = 4'b0001;
	ROM[830] = 4'b0000;
	ROM[831] = 4'b0000;
	ROM[832] = 4'b0000;
	ROM[833] = 4'b0100;
	ROM[834] = 4'b0000;
	ROM[835] = 4'b0100;
	ROM[836] = 4'b0000;
	ROM[837] = 4'b0100;
	ROM[838] = 4'b0000;
	ROM[839] = 4'b0000;
	ROM[840] = 4'b0000;
	ROM[841] = 4'b0001;
	ROM[842] = 4'b0000;
	ROM[843] = 4'b0001;
	ROM[844] = 4'b0000;
	ROM[845] = 4'b0001;
	ROM[846] = 4'b0000;
	ROM[847] = 4'b0000;
	ROM[848] = 4'b0000;
	ROM[849] = 4'b0100;
	ROM[850] = 4'b0000;
	ROM[851] = 4'b0000;
	ROM[852] = 4'b0000;
	ROM[853] = 4'b0010;
	ROM[854] = 4'b0011;
	ROM[855] = 4'b0011;
	ROM[856] = 4'b0011;
	ROM[857] = 4'b1011;
	ROM[858] = 4'b1100;
	ROM[859] = 4'b1100;
	ROM[860] = 4'b1100;
	ROM[861] = 4'b1101;
	ROM[862] = 4'b0000;
	ROM[863] = 4'b0000;
	ROM[864] = 4'b0000;
	ROM[865] = 4'b0101;
	ROM[866] = 4'b0000;
	ROM[867] = 4'b0000;
	ROM[868] = 4'b0000;
	ROM[869] = 4'b0100;
	ROM[870] = 4'b0000;
	ROM[871] = 4'b0000;
	ROM[872] = 4'b0000;
	ROM[873] = 4'b0000;
	ROM[874] = 4'b0000;
	ROM[875] = 4'b0000;
	ROM[876] = 4'b0000;
	ROM[877] = 4'b0100;
	ROM[878] = 4'b0000;
	ROM[879] = 4'b0000;
	ROM[880] = 4'b0000;
	ROM[881] = 4'b0000;
	ROM[882] = 4'b0000;
	ROM[883] = 4'b0000;
	ROM[884] = 4'b0000;
	ROM[885] = 4'b0100;
	ROM[886] = 4'b0000;
	ROM[887] = 4'b0000;
	ROM[888] = 4'b0000;
	ROM[889] = 4'b0000;
	ROM[890] = 4'b0000;
	ROM[891] = 4'b0000;
	ROM[892] = 4'b0000;
	ROM[893] = 4'b0100;
	ROM[894] = 4'b0000;
	ROM[895] = 4'b0000;
	ROM[896] = 4'b0000;
	ROM[897] = 4'b0001;
	ROM[898] = 4'b0000;
	ROM[899] = 4'b0000;
	ROM[900] = 4'b0000;
	ROM[901] = 4'b0100;
	ROM[902] = 4'b0000;
	ROM[903] = 4'b0000;
	ROM[904] = 4'b0000;
	ROM[905] = 4'b0001;
	ROM[906] = 4'b0000;
	ROM[907] = 4'b0000;
	ROM[908] = 4'b0000;
	ROM[909] = 4'b0100;
	ROM[910] = 4'b0000;
	ROM[911] = 4'b0000;
	ROM[912] = 4'b0000;
	ROM[913] = 4'b1000;
	ROM[914] = 4'b1100;
	ROM[915] = 4'b1100;
	ROM[916] = 4'b1100;
	ROM[917] = 4'b1100;
	ROM[918] = 4'b1100;
	ROM[919] = 4'b1100;
	ROM[920] = 4'b1100;
	ROM[921] = 4'b1100;
	ROM[922] = 4'b1100;
	ROM[923] = 4'b1100;
	ROM[924] = 4'b1100;
	ROM[925] = 4'b1100;
	ROM[926] = 4'b1100;
	ROM[927] = 4'b1100;
	ROM[928] = 4'b1100;
	ROM[929] = 4'b1110;
	ROM[930] = 4'b0011;
	ROM[931] = 4'b0011;
	ROM[932] = 4'b0011;
	ROM[933] = 4'b0111;
	ROM[934] = 4'b0000;
	ROM[935] = 4'b0100;
	ROM[936] = 4'b0000;
	ROM[937] = 4'b0001;
	ROM[938] = 4'b0000;
	ROM[939] = 4'b0001;
	ROM[940] = 4'b0000;
	ROM[941] = 4'b0100;
	ROM[942] = 4'b0000;
	ROM[943] = 4'b0100;
	ROM[944] = 4'b0000;
	ROM[945] = 4'b0001;
	ROM[946] = 4'b0000;
	ROM[947] = 4'b0001;
	ROM[948] = 4'b0000;
	ROM[949] = 4'b0100;
	ROM[950] = 4'b0000;
	ROM[951] = 4'b0100;
	ROM[952] = 4'b0000;
	ROM[953] = 4'b0001;
	ROM[954] = 4'b0000;
	ROM[955] = 4'b0010;
	ROM[956] = 4'b0011;
	ROM[957] = 4'b0011;
	ROM[958] = 4'b0011;
	ROM[959] = 4'b0111;
	ROM[960] = 4'b0000;
	ROM[961] = 4'b0100;
	ROM[962] = 4'b0000;
	ROM[963] = 4'b0001;
	ROM[964] = 4'b0000;
	ROM[965] = 4'b0010;
	ROM[966] = 4'b0011;
	ROM[967] = 4'b0011;
	ROM[968] = 4'b0011;
	ROM[969] = 4'b0111;
	ROM[970] = 4'b0000;
	ROM[971] = 4'b0100;
	ROM[972] = 4'b0000;
	ROM[973] = 4'b0001;
	ROM[974] = 4'b0000;
	ROM[975] = 4'b0001;
	ROM[976] = 4'b0000;
	ROM[977] = 4'b0100;
	ROM[978] = 4'b0000;
	ROM[979] = 4'b0100;
	ROM[980] = 4'b0000;
	ROM[981] = 4'b0001;
	ROM[982] = 4'b0000;
	ROM[983] = 4'b0001;
	ROM[984] = 4'b0000;
	ROM[985] = 4'b0010;
	ROM[986] = 4'b0011;
	ROM[987] = 4'b0011;
	ROM[988] = 4'b0011;
	ROM[989] = 4'b0011;
	ROM[990] = 4'b0011;
	ROM[991] = 4'b0011;
	ROM[992] = 4'b0011;
	ROM[993] = 4'b1011;
	ROM[994] = 4'b1100;
	ROM[995] = 4'b1100;
	ROM[996] = 4'b1100;
	ROM[997] = 4'b1101;
	ROM[998] = 4'b0000;
	ROM[999] = 4'b0001;
	ROM[1000] = 4'b0000;
	ROM[1001] = 4'b0100;
	ROM[1002] = 4'b0000;
	ROM[1003] = 4'b0100;
	ROM[1004] = 4'b0000;
	ROM[1005] = 4'b0001;
	ROM[1006] = 4'b0000;
	ROM[1007] = 4'b0001;
	ROM[1008] = 4'b0000;
	ROM[1009] = 4'b0100;
	ROM[1010] = 4'b0000;
	ROM[1011] = 4'b0100;
	ROM[1012] = 4'b0000;
	ROM[1013] = 4'b0001;
	ROM[1014] = 4'b0000;
	ROM[1015] = 4'b0001;
	ROM[1016] = 4'b0000;
	ROM[1017] = 4'b0100;
	ROM[1018] = 4'b0000;
	ROM[1019] = 4'b1000;
	ROM[1020] = 4'b1100;
	ROM[1021] = 4'b1100;
	ROM[1022] = 4'b1100;
	ROM[1023] = 4'b1101;
	ROM[1024] = 4'b0000;
	ROM[1025] = 4'b0100;
	ROM[1026] = 4'b0000;
	ROM[1027] = 4'b0100;
	ROM[1028] = 4'b0000;
	ROM[1029] = 4'b0100;
	ROM[1030] = 4'b0000;
	ROM[1031] = 4'b0100;
	ROM[1032] = 4'b0000;
	ROM[1033] = 4'b0001;
	ROM[1034] = 4'b0000;
	ROM[1035] = 4'b0001;
	ROM[1036] = 4'b0000;
	ROM[1037] = 4'b0001;
	ROM[1038] = 4'b0000;
	ROM[1039] = 4'b0001;
	ROM[1040] = 4'b0000;
	ROM[1041] = 4'b0100;
	ROM[1042] = 4'b0000;
	ROM[1043] = 4'b0000;
	ROM[1044] = 4'b0100;
	ROM[1045] = 4'b0000;
	ROM[1046] = 4'b0000;
	ROM[1047] = 4'b0001;
	ROM[1048] = 4'b0000;
	ROM[1049] = 4'b0001;
	ROM[1050] = 4'b0000;
	ROM[1051] = 4'b0000;
	ROM[1052] = 4'b0000;
	ROM[1053] = 4'b0100;
	ROM[1054] = 4'b0000;
	ROM[1055] = 4'b0000;
	ROM[1056] = 4'b0000;
	ROM[1057] = 4'b0010;
	ROM[1058] = 4'b0011;
	ROM[1059] = 4'b0011;
	ROM[1060] = 4'b0011;
	ROM[1061] = 4'b0111;
	ROM[1062] = 4'b0000;
	ROM[1063] = 4'b0100;
	ROM[1064] = 4'b0000;
	ROM[1065] = 4'b0001;
	ROM[1066] = 4'b0000;
	ROM[1067] = 4'b0001;
	ROM[1068] = 4'b0000;
	ROM[1069] = 4'b0100;
	ROM[1070] = 4'b0000;
	ROM[1071] = 4'b0100;
	ROM[1072] = 4'b0000;
	ROM[1073] = 4'b0001;
	ROM[1074] = 4'b0000;
	ROM[1075] = 4'b0001;
	ROM[1076] = 4'b0000;
	ROM[1077] = 4'b0100;
	ROM[1078] = 4'b0000;
	ROM[1079] = 4'b0100;
	ROM[1080] = 4'b0000;
	ROM[1081] = 4'b0001;
	ROM[1082] = 4'b0000;
	ROM[1083] = 4'b0010;
	ROM[1084] = 4'b0011;
	ROM[1085] = 4'b0011;
	ROM[1086] = 4'b0011;
	ROM[1087] = 4'b0111;
	ROM[1088] = 4'b0000;
	ROM[1089] = 4'b0100;
	ROM[1090] = 4'b0000;
	ROM[1091] = 4'b0001;
	ROM[1092] = 4'b0000;
	ROM[1093] = 4'b0010;
	ROM[1094] = 4'b0011;
	ROM[1095] = 4'b0011;
	ROM[1096] = 4'b0011;
	ROM[1097] = 4'b0111;
	ROM[1098] = 4'b0000;
	ROM[1099] = 4'b0100;
	ROM[1100] = 4'b0000;
	ROM[1101] = 4'b0001;
	ROM[1102] = 4'b0000;
	ROM[1103] = 4'b0001;
	ROM[1104] = 4'b0000;
	ROM[1105] = 4'b1000;
	ROM[1106] = 4'b1100;
	ROM[1107] = 4'b1100;
	ROM[1108] = 4'b1100;
	ROM[1109] = 4'b1100;
	ROM[1110] = 4'b1100;
	ROM[1111] = 4'b1100;
	ROM[1112] = 4'b1100;
	ROM[1113] = 4'b1110;
	ROM[1114] = 4'b0011;
	ROM[1115] = 4'b0011;
	ROM[1116] = 4'b0011;
	ROM[1117] = 4'b0011;
	ROM[1118] = 4'b0011;
	ROM[1119] = 4'b0011;
	ROM[1120] = 4'b0011;
	ROM[1121] = 4'b0111;
	ROM[1122] = 4'b0000;
	ROM[1123] = 4'b0100;
	ROM[1124] = 4'b0000;
	ROM[1125] = 4'b0100;
	ROM[1126] = 4'b0000;
	ROM[1127] = 4'b0100;
	ROM[1128] = 4'b0000;
	ROM[1129] = 4'b0001;
	ROM[1130] = 4'b0000;
	ROM[1131] = 4'b0001;
	ROM[1132] = 4'b0000;
	ROM[1133] = 4'b0001;
	ROM[1134] = 4'b0000;
	ROM[1135] = 4'b0001;
	ROM[1136] = 4'b0000;
	ROM[1137] = 4'b0100;
	ROM[1138] = 4'b0000;
	ROM[1139] = 4'b0000;
	ROM[1140] = 4'b0100;
	ROM[1141] = 4'b0000;
	ROM[1142] = 4'b0000;
	ROM[1143] = 4'b0001;
	ROM[1144] = 4'b0000;
	ROM[1145] = 4'b0001;
	ROM[1146] = 4'b0000;
	ROM[1147] = 4'b0000;
	ROM[1148] = 4'b0000;
	ROM[1149] = 4'b0100;
	ROM[1150] = 4'b0000;
	ROM[1151] = 4'b0000;
	ROM[1152] = 4'b0000;
	ROM[1153] = 4'b0001;
	ROM[1154] = 4'b0000;
	ROM[1155] = 4'b0001;
	ROM[1156] = 4'b0000;
	ROM[1157] = 4'b0001;
	ROM[1158] = 4'b0000;
	ROM[1159] = 4'b0001;
	ROM[1160] = 4'b0000;
	ROM[1161] = 4'b0100;
	ROM[1162] = 4'b0000;
	ROM[1163] = 4'b0100;
	ROM[1164] = 4'b0000;
	ROM[1165] = 4'b0100;
	ROM[1166] = 4'b0000;
	ROM[1167] = 4'b0100;
	ROM[1168] = 4'b0000;
	ROM[1169] = 4'b0010;
	ROM[1170] = 4'b0011;
	ROM[1171] = 4'b0011;
	ROM[1172] = 4'b0011;
	ROM[1173] = 4'b0011;
	ROM[1174] = 4'b0011;
	ROM[1175] = 4'b0011;
	ROM[1176] = 4'b0011;
	ROM[1177] = 4'b0011;
	ROM[1178] = 4'b0011;
	ROM[1179] = 4'b0011;
	ROM[1180] = 4'b0011;
	ROM[1181] = 4'b0011;
	ROM[1182] = 4'b0011;
	ROM[1183] = 4'b0011;
	ROM[1184] = 4'b0011;
	ROM[1185] = 4'b0111;
	ROM[1186] = 4'b0000;
	ROM[1187] = 4'b0000;
	ROM[1188] = 4'b0000;
	ROM[1189] = 4'b0000;
	ROM[1190] = 4'b0000;
	ROM[1191] = 4'b0100;
	ROM[1192] = 4'b0000;
	ROM[1193] = 4'b0000;
	ROM[1194] = 4'b0000;
	ROM[1195] = 4'b0000;
	ROM[1196] = 4'b0000;
	ROM[1197] = 4'b0001;
	ROM[1198] = 4'b0000;
	ROM[1199] = 4'b0000;
	ROM[1200] = 4'b0000;
	ROM[1201] = 4'b0000;
	ROM[1202] = 4'b0000;
	ROM[1203] = 4'b0100;
	ROM[1204] = 4'b0000;
	ROM[1205] = 4'b0100;
	ROM[1206] = 4'b0000;
	ROM[1207] = 4'b0000;
	ROM[1208] = 4'b0000;
	ROM[1209] = 4'b0001;
	ROM[1210] = 4'b0000;
	ROM[1211] = 4'b0000;
	ROM[1212] = 4'b0000;
	ROM[1213] = 4'b0100;
	ROM[1214] = 4'b0000;
	ROM[1215] = 4'b0000;
	ROM[1216] = 4'b0000;
	ROM[1217] = 4'b0001;
	ROM[1218] = 4'b0000;
	ROM[1219] = 4'b0000;
	ROM[1220] = 4'b0000;
	ROM[1221] = 4'b0100;
	ROM[1222] = 4'b0000;
	ROM[1223] = 4'b0000;
	ROM[1224] = 4'b0000;
	ROM[1225] = 4'b0001;
	ROM[1226] = 4'b0000;
	ROM[1227] = 4'b0001;
	ROM[1228] = 4'b0000;
	ROM[1229] = 4'b0000;
	ROM[1230] = 4'b0000;
	ROM[1231] = 4'b0100;
	ROM[1232] = 4'b0000;
	ROM[1233] = 4'b0100;
	ROM[1234] = 4'b0000;
	ROM[1235] = 4'b0100;
	ROM[1236] = 4'b0000;
	ROM[1237] = 4'b0000;
	ROM[1238] = 4'b0000;
	ROM[1239] = 4'b0000;
	ROM[1240] = 4'b0000;
	ROM[1241] = 4'b0000;
	ROM[1242] = 4'b0000;
	ROM[1243] = 4'b0001;
	ROM[1244] = 4'b0000;
	ROM[1245] = 4'b0000;
	ROM[1246] = 4'b0000;
	ROM[1247] = 4'b0000;
	ROM[1248] = 4'b0000;
	ROM[1249] = 4'b0100;
	ROM[1250] = 4'b0000;
	ROM[1251] = 4'b0000;
	ROM[1252] = 4'b0000;
	ROM[1253] = 4'b0000;
	ROM[1254] = 4'b0000;
	ROM[1255] = 4'b0001;
	ROM[1256] = 4'b0000;
	ROM[1257] = 4'b0000;
	ROM[1258] = 4'b0000;
	ROM[1259] = 4'b0000;
	ROM[1260] = 4'b0000;
	ROM[1261] = 4'b0100;
	ROM[1262] = 4'b0000;
	ROM[1263] = 4'b0000;
	ROM[1264] = 4'b0000;
	ROM[1265] = 4'b0000;
	ROM[1266] = 4'b0000;
	ROM[1267] = 4'b0001;
	ROM[1268] = 4'b0000;
	ROM[1269] = 4'b0001;
	ROM[1270] = 4'b0000;
	ROM[1271] = 4'b0000;
	ROM[1272] = 4'b0000;
	ROM[1273] = 4'b0100;
	ROM[1274] = 4'b0000;
	ROM[1275] = 4'b0000;
	ROM[1276] = 4'b0000;
	ROM[1277] = 4'b0001;
	ROM[1278] = 4'b0000;
	ROM[1279] = 4'b0000;
	ROM[1280] = 4'b0000;
	ROM[1281] = 4'b0100;
	ROM[1282] = 4'b0000;
	ROM[1283] = 4'b0000;
	ROM[1284] = 4'b0000;
	ROM[1285] = 4'b0001;
	ROM[1286] = 4'b0000;
	ROM[1287] = 4'b0000;
	ROM[1288] = 4'b0000;
	ROM[1289] = 4'b0100;
	ROM[1290] = 4'b0000;
	ROM[1291] = 4'b0100;
	ROM[1292] = 4'b0000;
	ROM[1293] = 4'b0000;
	ROM[1294] = 4'b0000;
	ROM[1295] = 4'b0001;
	ROM[1296] = 4'b0000;
	ROM[1297] = 4'b0001;
	ROM[1298] = 4'b0000;
	ROM[1299] = 4'b0001;
	ROM[1300] = 4'b0000;
	ROM[1301] = 4'b0000;
	ROM[1302] = 4'b0000;
	ROM[1303] = 4'b0000;
	ROM[1304] = 4'b0000;
	ROM[1305] = 4'b1000;
	ROM[1306] = 4'b1100;
	ROM[1307] = 4'b1100;
	ROM[1308] = 4'b1100;
	ROM[1309] = 4'b1101;
	ROM[1310] = 4'b0000;
	ROM[1311] = 4'b0000;
	ROM[1312] = 4'b0000;
	ROM[1313] = 4'b0101;
	ROM[1314] = 4'b0000;
	ROM[1315] = 4'b0000;
	ROM[1316] = 4'b0000;
	ROM[1317] = 4'b0000;
	ROM[1318] = 4'b0000;
	ROM[1319] = 4'b0100;
	ROM[1320] = 4'b0000;
	ROM[1321] = 4'b0000;
	ROM[1322] = 4'b0000;
	ROM[1323] = 4'b0001;
	ROM[1324] = 4'b0000;
	ROM[1325] = 4'b0001;
	ROM[1326] = 4'b0000;
	ROM[1327] = 4'b0000;
	ROM[1328] = 4'b0000;
	ROM[1329] = 4'b0100;
	ROM[1330] = 4'b0000;
	ROM[1331] = 4'b0000;
	ROM[1332] = 4'b0000;
	ROM[1333] = 4'b0001;
	ROM[1334] = 4'b0000;
	ROM[1335] = 4'b0000;
	ROM[1336] = 4'b0000;
	ROM[1337] = 4'b0100;
	ROM[1338] = 4'b0000;
	ROM[1339] = 4'b0000;
	ROM[1340] = 4'b0000;
	ROM[1341] = 4'b0001;
	ROM[1342] = 4'b0000;
	ROM[1343] = 4'b0000;
	ROM[1344] = 4'b0000;
	ROM[1345] = 4'b0100;
	ROM[1346] = 4'b0000;
	ROM[1347] = 4'b0000;
	ROM[1348] = 4'b0000;
	ROM[1349] = 4'b0001;
	ROM[1350] = 4'b0000;
	ROM[1351] = 4'b0000;
	ROM[1352] = 4'b0000;
	ROM[1353] = 4'b0100;
	ROM[1354] = 4'b0000;
	ROM[1355] = 4'b0100;
	ROM[1356] = 4'b0000;
	ROM[1357] = 4'b0000;
	ROM[1358] = 4'b0000;
	ROM[1359] = 4'b0001;
	ROM[1360] = 4'b0000;
	ROM[1361] = 4'b0001;
	ROM[1362] = 4'b0000;
	ROM[1363] = 4'b0001;
	ROM[1364] = 4'b0000;
	ROM[1365] = 4'b0000;
	ROM[1366] = 4'b0000;
	ROM[1367] = 4'b0000;
	ROM[1368] = 4'b0000;
	ROM[1369] = 4'b0000;
	ROM[1370] = 4'b0000;
	ROM[1371] = 4'b0100;
	ROM[1372] = 4'b0000;
	ROM[1373] = 4'b0000;
	ROM[1374] = 4'b0000;
	ROM[1375] = 4'b0000;
	ROM[1376] = 4'b0000;
	ROM[1377] = 4'b0101;
	ROM[1378] = 4'b0000;
	ROM[1379] = 4'b0000;
	ROM[1380] = 4'b0000;
	ROM[1381] = 4'b0000;
	ROM[1382] = 4'b0000;
	ROM[1383] = 4'b0001;
	ROM[1384] = 4'b0000;
	ROM[1385] = 4'b0000;
	ROM[1386] = 4'b0000;
	ROM[1387] = 4'b0100;
	ROM[1388] = 4'b0000;
	ROM[1389] = 4'b0100;
	ROM[1390] = 4'b0000;
	ROM[1391] = 4'b0000;
	ROM[1392] = 4'b0000;
	ROM[1393] = 4'b0001;
	ROM[1394] = 4'b0000;
	ROM[1395] = 4'b0000;
	ROM[1396] = 4'b0000;
	ROM[1397] = 4'b0100;
	ROM[1398] = 4'b0000;
	ROM[1399] = 4'b0000;
	ROM[1400] = 4'b0000;
	ROM[1401] = 4'b0001;
	ROM[1402] = 4'b0000;
	ROM[1403] = 4'b0000;
	ROM[1404] = 4'b0000;
	ROM[1405] = 4'b0100;
	ROM[1406] = 4'b0000;
	ROM[1407] = 4'b0000;
	ROM[1408] = 4'b0000;
	ROM[1409] = 4'b0001;
	ROM[1410] = 4'b0000;
	ROM[1411] = 4'b0000;
	ROM[1412] = 4'b0000;
	ROM[1413] = 4'b0100;
	ROM[1414] = 4'b0000;
	ROM[1415] = 4'b0000;
	ROM[1416] = 4'b0000;
	ROM[1417] = 4'b0001;
	ROM[1418] = 4'b0000;
	ROM[1419] = 4'b0001;
	ROM[1420] = 4'b0000;
	ROM[1421] = 4'b0000;
	ROM[1422] = 4'b0000;
	ROM[1423] = 4'b0100;
	ROM[1424] = 4'b0000;
	ROM[1425] = 4'b1000;
	ROM[1426] = 4'b1100;
	ROM[1427] = 4'b1100;
	ROM[1428] = 4'b1100;
	ROM[1429] = 4'b1100;
	ROM[1430] = 4'b1100;
	ROM[1431] = 4'b1100;
	ROM[1432] = 4'b1100;
	ROM[1433] = 4'b1100;
	ROM[1434] = 4'b1100;
	ROM[1435] = 4'b1100;
	ROM[1436] = 4'b1100;
	ROM[1437] = 4'b1100;
	ROM[1438] = 4'b1100;
	ROM[1439] = 4'b1100;
	ROM[1440] = 4'b1100;
	ROM[1441] = 4'b1101;
	ROM[1442] = 4'b0000;
	ROM[1443] = 4'b0000;
	ROM[1444] = 4'b0000;
	ROM[1445] = 4'b0001;
	ROM[1446] = 4'b0000;
	ROM[1447] = 4'b0000;
	ROM[1448] = 4'b0000;
	ROM[1449] = 4'b0001;
	ROM[1450] = 4'b0000;
	ROM[1451] = 4'b0000;
	ROM[1452] = 4'b0000;
	ROM[1453] = 4'b0100;
	ROM[1454] = 4'b0000;
	ROM[1455] = 4'b0100;
	ROM[1456] = 4'b0000;
	ROM[1457] = 4'b0100;
	ROM[1458] = 4'b0000;
	ROM[1459] = 4'b0000;
	ROM[1460] = 4'b0000;
	ROM[1461] = 4'b0100;
	ROM[1462] = 4'b0000;
	ROM[1463] = 4'b0000;
	ROM[1464] = 4'b0000;
	ROM[1465] = 4'b0001;
	ROM[1466] = 4'b0000;
	ROM[1467] = 4'b0001;
	ROM[1468] = 4'b0000;
	ROM[1469] = 4'b0001;
	ROM[1470] = 4'b0000;
	ROM[1471] = 4'b0001;
	ROM[1472] = 4'b0000;
	ROM[1473] = 4'b0100;
	ROM[1474] = 4'b0000;
	ROM[1475] = 4'b0100;
	ROM[1476] = 4'b0000;
	ROM[1477] = 4'b0100;
	ROM[1478] = 4'b0000;
	ROM[1479] = 4'b0000;
	ROM[1480] = 4'b0000;
	ROM[1481] = 4'b0100;
	ROM[1482] = 4'b0000;
	ROM[1483] = 4'b0000;
	ROM[1484] = 4'b0000;
	ROM[1485] = 4'b0001;
	ROM[1486] = 4'b0000;
	ROM[1487] = 4'b0001;
	ROM[1488] = 4'b0000;
	ROM[1489] = 4'b0001;
	ROM[1490] = 4'b0000;
	ROM[1491] = 4'b0000;
	ROM[1492] = 4'b0000;
	ROM[1493] = 4'b0001;
	ROM[1494] = 4'b0000;
	ROM[1495] = 4'b0000;
	ROM[1496] = 4'b0000;
	ROM[1497] = 4'b0100;
	ROM[1498] = 4'b0000;
	ROM[1499] = 4'b0100;
	ROM[1500] = 4'b0000;
	ROM[1501] = 4'b0100;
	ROM[1502] = 4'b0000;
	ROM[1503] = 4'b0100;
	ROM[1504] = 4'b0000;
	ROM[1505] = 4'b0001;
	ROM[1506] = 4'b0000;
	ROM[1507] = 4'b0001;
	ROM[1508] = 4'b0000;
	ROM[1509] = 4'b0001;
	ROM[1510] = 4'b0000;
	ROM[1511] = 4'b0000;
	ROM[1512] = 4'b0000;
	ROM[1513] = 4'b0001;
	ROM[1514] = 4'b0000;
	ROM[1515] = 4'b0000;
	ROM[1516] = 4'b0000;
	ROM[1517] = 4'b0100;
	ROM[1518] = 4'b0000;
	ROM[1519] = 4'b0100;
	ROM[1520] = 4'b0000;
	ROM[1521] = 4'b0100;
	ROM[1522] = 4'b0000;
	ROM[1523] = 4'b0000;
	ROM[1524] = 4'b0000;
	ROM[1525] = 4'b0100;
	ROM[1526] = 4'b0000;
	ROM[1527] = 4'b0000;
	ROM[1528] = 4'b0000;
	ROM[1529] = 4'b0001;
	ROM[1530] = 4'b0000;
	ROM[1531] = 4'b0001;
	ROM[1532] = 4'b0000;
	ROM[1533] = 4'b0001;
	ROM[1534] = 4'b0000;
	ROM[1535] = 4'b0001;
	ROM[1536] = 4'b0000;
	ROM[1537] = 4'b0100;
	ROM[1538] = 4'b0000;
	ROM[1539] = 4'b0100;
	ROM[1540] = 4'b0000;
	ROM[1541] = 4'b0100;
	ROM[1542] = 4'b0000;
	ROM[1543] = 4'b0100;
	ROM[1544] = 4'b0000;
	ROM[1545] = 4'b0001;
	ROM[1546] = 4'b0000;
	ROM[1547] = 4'b0001;
	ROM[1548] = 4'b0000;
	ROM[1549] = 4'b0001;
	ROM[1550] = 4'b0000;
	ROM[1551] = 4'b0001;
	ROM[1552] = 4'b0000;
	ROM[1553] = 4'b1000;
	ROM[1554] = 4'b1100;
	ROM[1555] = 4'b1100;
	ROM[1556] = 4'b1100;
	ROM[1557] = 4'b1100;
	ROM[1558] = 4'b1100;
	ROM[1559] = 4'b1100;
	ROM[1560] = 4'b1100;
	ROM[1561] = 4'b1100;
	ROM[1562] = 4'b1100;
	ROM[1563] = 4'b1100;
	ROM[1564] = 4'b1100;
	ROM[1565] = 4'b1100;
	ROM[1566] = 4'b1100;
	ROM[1567] = 4'b1100;
	ROM[1568] = 4'b1100;
	ROM[1569] = 4'b1100;
	ROM[1570] = 4'b0000;
	ROM[1571] = 4'b0000;
	ROM[1572] = 4'b0000;
	ROM[1573] = 4'b0000;
	ROM[1574] = 4'b0000;
	ROM[1575] = 4'b0000;
	ROM[1576] = 4'b0000;
	ROM[1577] = 4'b0000;
	ROM[1578] = 4'b0000;
	ROM[1579] = 4'b0000;
	ROM[1580] = 4'b0000;
	ROM[1581] = 4'b0000;
	ROM[1582] = 4'b0000;
	ROM[1583] = 4'b0000;
	ROM[1584] = 4'b0000;
	ROM[1585] = 4'b0100;
	ROM[1586] = 4'b0000;
	ROM[1587] = 4'b0000;
	ROM[1588] = 4'b0000;
	ROM[1589] = 4'b0000;
	ROM[1590] = 4'b0000;
	ROM[1591] = 4'b0000;
	ROM[1592] = 4'b0000;
	ROM[1593] = 4'b0000;
	ROM[1594] = 4'b0000;
	ROM[1595] = 4'b0000;
	ROM[1596] = 4'b0000;
	ROM[1597] = 4'b0001;
	ROM[1598] = 4'b0000;
	ROM[1599] = 4'b0000;
	ROM[1600] = 4'b0000;
	ROM[1601] = 4'b0010;
	ROM[1602] = 4'b0011;
	ROM[1603] = 4'b0011;
	ROM[1604] = 4'b0000;
	ROM[1605] = 4'b0100;
	ROM[1606] = 4'b0000;
	ROM[1607] = 4'b1000;
	ROM[1608] = 4'b1100;
	ROM[1609] = 4'b1100;
	ROM[1610] = 4'b0000;
	ROM[1611] = 4'b0010;
	ROM[1612] = 4'b0011;
	ROM[1613] = 4'b0011;
	ROM[1614] = 4'b0000;
	ROM[1615] = 4'b0100;
	ROM[1616] = 4'b0000;
	ROM[1617] = 4'b1000;
	ROM[1618] = 4'b1100;
	ROM[1619] = 4'b1100;
	ROM[1620] = 4'b0000;
	ROM[1621] = 4'b0001;
	ROM[1622] = 4'b0000;
	ROM[1623] = 4'b0010;
	ROM[1624] = 4'b0011;
	ROM[1625] = 4'b0011;
	ROM[1626] = 4'b0000;
	ROM[1627] = 4'b1000;
	ROM[1628] = 4'b1100;
	ROM[1629] = 4'b1100;
	ROM[1630] = 4'b0000;
	ROM[1631] = 4'b0001;
	ROM[1632] = 4'b0000;
	ROM[1633] = 4'b0010;
	ROM[1634] = 4'b0011;
	ROM[1635] = 4'b0011;
	ROM[1636] = 4'b0000;
	ROM[1637] = 4'b0100;
	ROM[1638] = 4'b0000;
	ROM[1639] = 4'b0100;
	ROM[1640] = 4'b0000;
	ROM[1641] = 4'b1000;
	ROM[1642] = 4'b1100;
	ROM[1643] = 4'b1100;
	ROM[1644] = 4'b0000;
	ROM[1645] = 4'b0001;
	ROM[1646] = 4'b0000;
	ROM[1647] = 4'b0001;
	ROM[1648] = 4'b0000;
	ROM[1649] = 4'b0100;
	ROM[1650] = 4'b0000;
	ROM[1651] = 4'b0100;
	ROM[1652] = 4'b0000;
	ROM[1653] = 4'b0001;
	ROM[1654] = 4'b0000;
	ROM[1655] = 4'b0001;
	ROM[1656] = 4'b0000;
	ROM[1657] = 4'b0000;
	ROM[1658] = 4'b0000;
	ROM[1659] = 4'b0100;
	ROM[1660] = 4'b0000;
	ROM[1661] = 4'b0100;
	ROM[1662] = 4'b0000;
	ROM[1663] = 4'b0001;
	ROM[1664] = 4'b0000;
	ROM[1665] = 4'b0010;
	ROM[1666] = 4'b0011;
	ROM[1667] = 4'b0011;
	ROM[1668] = 4'b0000;
	ROM[1669] = 4'b0100;
	ROM[1670] = 4'b0000;
	ROM[1671] = 4'b1000;
	ROM[1672] = 4'b1100;
	ROM[1673] = 4'b1100;
	ROM[1674] = 4'b0000;
	ROM[1675] = 4'b0010;
	ROM[1676] = 4'b0011;
	ROM[1677] = 4'b0011;
	ROM[1678] = 4'b0000;
	ROM[1679] = 4'b0100;
	ROM[1680] = 4'b0000;
	ROM[1681] = 4'b1000;
	ROM[1682] = 4'b1100;
	ROM[1683] = 4'b1100;
	ROM[1684] = 4'b0000;
	ROM[1685] = 4'b0001;
	ROM[1686] = 4'b0000;
	ROM[1687] = 4'b0010;
	ROM[1688] = 4'b0011;
	ROM[1689] = 4'b0011;
	ROM[1690] = 4'b0000;
	ROM[1691] = 4'b1000;
	ROM[1692] = 4'b1100;
	ROM[1693] = 4'b1100;
	ROM[1694] = 4'b0000;
	ROM[1695] = 4'b0001;
	ROM[1696] = 4'b0000;
	ROM[1697] = 4'b0100;
	ROM[1698] = 4'b0000;
	ROM[1699] = 4'b0100;
	ROM[1700] = 4'b0000;
	ROM[1701] = 4'b0001;
	ROM[1702] = 4'b0000;
	ROM[1703] = 4'b0001;
	ROM[1704] = 4'b0000;
	ROM[1705] = 4'b0100;
	ROM[1706] = 4'b0000;
	ROM[1707] = 4'b0100;
	ROM[1708] = 4'b0000;
	ROM[1709] = 4'b0001;
	ROM[1710] = 4'b0000;
	ROM[1711] = 4'b0001;
	ROM[1712] = 4'b0000;
	ROM[1713] = 4'b0100;
	ROM[1714] = 4'b0000;
	ROM[1715] = 4'b0000;
	ROM[1716] = 4'b0100;
	ROM[1717] = 4'b0000;
	ROM[1718] = 4'b0000;
	ROM[1719] = 4'b0001;
	ROM[1720] = 4'b0000;
	ROM[1721] = 4'b0001;
	ROM[1722] = 4'b0000;
	ROM[1723] = 4'b0000;
	ROM[1724] = 4'b0000;
	ROM[1725] = 4'b0100;
	ROM[1726] = 4'b0000;
	ROM[1727] = 4'b0000;
	ROM[1728] = 4'b0000;
	ROM[1729] = 4'b1000;
	ROM[1730] = 4'b1100;
	ROM[1731] = 4'b1100;
	ROM[1732] = 4'b0000;
	ROM[1733] = 4'b0001;
	ROM[1734] = 4'b0000;
	ROM[1735] = 4'b0010;
	ROM[1736] = 4'b0011;
	ROM[1737] = 4'b0011;
	ROM[1738] = 4'b0000;
	ROM[1739] = 4'b1000;
	ROM[1740] = 4'b1100;
	ROM[1741] = 4'b1100;
	ROM[1742] = 4'b0000;
	ROM[1743] = 4'b0001;
	ROM[1744] = 4'b0000;
	ROM[1745] = 4'b0010;
	ROM[1746] = 4'b0011;
	ROM[1747] = 4'b0011;
	ROM[1748] = 4'b0000;
	ROM[1749] = 4'b0100;
	ROM[1750] = 4'b0000;
	ROM[1751] = 4'b1000;
	ROM[1752] = 4'b1100;
	ROM[1753] = 4'b1100;
	ROM[1754] = 4'b0000;
	ROM[1755] = 4'b0010;
	ROM[1756] = 4'b0011;
	ROM[1757] = 4'b0011;
	ROM[1758] = 4'b0000;
	ROM[1759] = 4'b0100;
	ROM[1760] = 4'b0000;
	ROM[1761] = 4'b1000;
	ROM[1762] = 4'b1100;
	ROM[1763] = 4'b1100;
	ROM[1764] = 4'b0000;
	ROM[1765] = 4'b0001;
	ROM[1766] = 4'b0000;
	ROM[1767] = 4'b0001;
	ROM[1768] = 4'b0000;
	ROM[1769] = 4'b0010;
	ROM[1770] = 4'b0011;
	ROM[1771] = 4'b0011;
	ROM[1772] = 4'b0000;
	ROM[1773] = 4'b0100;
	ROM[1774] = 4'b0000;
	ROM[1775] = 4'b0100;
	ROM[1776] = 4'b0000;
	ROM[1777] = 4'b0001;
	ROM[1778] = 4'b0000;
	ROM[1779] = 4'b0001;
	ROM[1780] = 4'b0000;
	ROM[1781] = 4'b0100;
	ROM[1782] = 4'b0000;
	ROM[1783] = 4'b0100;
	ROM[1784] = 4'b0000;
	ROM[1785] = 4'b0000;
	ROM[1786] = 4'b0000;
	ROM[1787] = 4'b0001;
	ROM[1788] = 4'b0000;
	ROM[1789] = 4'b0001;
	ROM[1790] = 4'b0000;
	ROM[1791] = 4'b0100;
	ROM[1792] = 4'b0000;
	ROM[1793] = 4'b1000;
	ROM[1794] = 4'b1100;
	ROM[1795] = 4'b1100;
	ROM[1796] = 4'b0000;
	ROM[1797] = 4'b0001;
	ROM[1798] = 4'b0000;
	ROM[1799] = 4'b0010;
	ROM[1800] = 4'b0011;
	ROM[1801] = 4'b0011;
	ROM[1802] = 4'b0000;
	ROM[1803] = 4'b1000;
	ROM[1804] = 4'b1100;
	ROM[1805] = 4'b1100;
	ROM[1806] = 4'b0000;
	ROM[1807] = 4'b0001;
	ROM[1808] = 4'b0000;
	ROM[1809] = 4'b0010;
	ROM[1810] = 4'b0011;
	ROM[1811] = 4'b0011;
	ROM[1812] = 4'b0000;
	ROM[1813] = 4'b0100;
	ROM[1814] = 4'b0000;
	ROM[1815] = 4'b1000;
	ROM[1816] = 4'b1100;
	ROM[1817] = 4'b1100;
	ROM[1818] = 4'b0000;
	ROM[1819] = 4'b0010;
	ROM[1820] = 4'b0011;
	ROM[1821] = 4'b0011;
	ROM[1822] = 4'b0000;
	ROM[1823] = 4'b0100;
	ROM[1824] = 4'b0000;
	ROM[1825] = 4'b0100;
	ROM[1826] = 4'b0000;
	ROM[1827] = 4'b0000;
	ROM[1828] = 4'b0000;
	ROM[1829] = 4'b0001;
	ROM[1830] = 4'b0000;
	ROM[1831] = 4'b0000;
	ROM[1832] = 4'b0000;
	ROM[1833] = 4'b0100;
	ROM[1834] = 4'b0000;
	ROM[1835] = 4'b0000;
	ROM[1836] = 4'b0000;
	ROM[1837] = 4'b0001;
	ROM[1838] = 4'b0000;
	ROM[1839] = 4'b0001;
	ROM[1840] = 4'b0000;
	ROM[1841] = 4'b0101;
	ROM[1842] = 4'b0000;
	ROM[1843] = 4'b0000;
	ROM[1844] = 4'b0000;
	ROM[1845] = 4'b0000;
	ROM[1846] = 4'b0000;
	ROM[1847] = 4'b0101;
	ROM[1848] = 4'b0000;
	ROM[1849] = 4'b0000;
	ROM[1850] = 4'b0000;
	ROM[1851] = 4'b0000;
	ROM[1852] = 4'b0000;
	ROM[1853] = 4'b0001;
	ROM[1854] = 4'b0000;
	ROM[1855] = 4'b0000;
	ROM[1856] = 4'b0000;
	ROM[1857] = 4'b1000;
	ROM[1858] = 4'b1100;
	ROM[1859] = 4'b1100;
	ROM[1860] = 4'b1100;
	ROM[1861] = 4'b1100;
	ROM[1862] = 4'b1100;
	ROM[1863] = 4'b1100;
	ROM[1864] = 4'b1100;
	ROM[1865] = 4'b1100;
	ROM[1866] = 4'b1100;
	ROM[1867] = 4'b1100;
	ROM[1868] = 4'b1100;
	ROM[1869] = 4'b1100;
	ROM[1870] = 4'b1100;
	ROM[1871] = 4'b1100;
	ROM[1872] = 4'b1100;
	ROM[1873] = 4'b1100;
	ROM[1874] = 4'b1100;
	ROM[1875] = 4'b1100;
	ROM[1876] = 4'b1100;
	ROM[1877] = 4'b1100;
	ROM[1878] = 4'b1100;
	ROM[1879] = 4'b1100;
	ROM[1880] = 4'b1100;
	ROM[1881] = 4'b1100;
	ROM[1882] = 4'b1100;
	ROM[1883] = 4'b1100;
	ROM[1884] = 4'b1100;
	ROM[1885] = 4'b1100;
	ROM[1886] = 4'b1100;
	ROM[1887] = 4'b1100;
	ROM[1888] = 4'b1100;
	ROM[1889] = 4'b1110;
	ROM[1890] = 4'b0011;
	ROM[1891] = 4'b0011;
	ROM[1892] = 4'b0000;
	ROM[1893] = 4'b1000;
	ROM[1894] = 4'b1100;
	ROM[1895] = 4'b1100;
	ROM[1896] = 4'b0000;
	ROM[1897] = 4'b0001;
	ROM[1898] = 4'b0000;
	ROM[1899] = 4'b0010;
	ROM[1900] = 4'b0011;
	ROM[1901] = 4'b0011;
	ROM[1902] = 4'b0000;
	ROM[1903] = 4'b0100;
	ROM[1904] = 4'b0000;
	ROM[1905] = 4'b1000;
	ROM[1906] = 4'b1100;
	ROM[1907] = 4'b1100;
	ROM[1908] = 4'b0000;
	ROM[1909] = 4'b0010;
	ROM[1910] = 4'b0011;
	ROM[1911] = 4'b0011;
	ROM[1912] = 4'b0000;
	ROM[1913] = 4'b0100;
	ROM[1914] = 4'b0000;
	ROM[1915] = 4'b0100;
	ROM[1916] = 4'b0000;
	ROM[1917] = 4'b0100;
	ROM[1918] = 4'b0000;
	ROM[1919] = 4'b0000;
	ROM[1920] = 4'b0000;
	ROM[1921] = 4'b0010;
	ROM[1922] = 4'b0011;
	ROM[1923] = 4'b0011;
	ROM[1924] = 4'b0000;
	ROM[1925] = 4'b0100;
	ROM[1926] = 4'b0000;
	ROM[1927] = 4'b1000;
	ROM[1928] = 4'b1100;
	ROM[1929] = 4'b1100;
	ROM[1930] = 4'b0000;
	ROM[1931] = 4'b0010;
	ROM[1932] = 4'b0011;
	ROM[1933] = 4'b0011;
	ROM[1934] = 4'b0000;
	ROM[1935] = 4'b0100;
	ROM[1936] = 4'b0000;
	ROM[1937] = 4'b1000;
	ROM[1938] = 4'b1100;
	ROM[1939] = 4'b1100;
	ROM[1940] = 4'b0000;
	ROM[1941] = 4'b0001;
	ROM[1942] = 4'b0000;
	ROM[1943] = 4'b0010;
	ROM[1944] = 4'b0011;
	ROM[1945] = 4'b0011;
	ROM[1946] = 4'b0000;
	ROM[1947] = 4'b1000;
	ROM[1948] = 4'b1100;
	ROM[1949] = 4'b1100;
	ROM[1950] = 4'b0000;
	ROM[1951] = 4'b0001;
	ROM[1952] = 4'b0000;
	ROM[1953] = 4'b0100;
	ROM[1954] = 4'b0000;
	ROM[1955] = 4'b0100;
	ROM[1956] = 4'b0000;
	ROM[1957] = 4'b0001;
	ROM[1958] = 4'b0000;
	ROM[1959] = 4'b0001;
	ROM[1960] = 4'b0000;
	ROM[1961] = 4'b0100;
	ROM[1962] = 4'b0000;
	ROM[1963] = 4'b0100;
	ROM[1964] = 4'b0000;
	ROM[1965] = 4'b0001;
	ROM[1966] = 4'b0000;
	ROM[1967] = 4'b0001;
	ROM[1968] = 4'b0000;
	ROM[1969] = 4'b0101;
	ROM[1970] = 4'b0000;
	ROM[1971] = 4'b0000;
	ROM[1972] = 4'b0000;
	ROM[1973] = 4'b0000;
	ROM[1974] = 4'b0000;
	ROM[1975] = 4'b0101;
	ROM[1976] = 4'b0000;
	ROM[1977] = 4'b0000;
	ROM[1978] = 4'b0000;
	ROM[1979] = 4'b0000;
	ROM[1980] = 4'b0000;
	ROM[1981] = 4'b0100;
	ROM[1982] = 4'b0000;
	ROM[1983] = 4'b0000;
	ROM[1984] = 4'b0000;
	ROM[1985] = 4'b1000;
	ROM[1986] = 4'b1100;
	ROM[1987] = 4'b1100;
	ROM[1988] = 4'b0000;
	ROM[1989] = 4'b0001;
	ROM[1990] = 4'b0000;
	ROM[1991] = 4'b0001;
	ROM[1992] = 4'b0000;
	ROM[1993] = 4'b0100;
	ROM[1994] = 4'b0000;
	ROM[1995] = 4'b0100;
	ROM[1996] = 4'b0000;
	ROM[1997] = 4'b0001;
	ROM[1998] = 4'b0000;
	ROM[1999] = 4'b0010;
	ROM[2000] = 4'b0011;
	ROM[2001] = 4'b0011;
	ROM[2002] = 4'b0000;
	ROM[2003] = 4'b0100;
	ROM[2004] = 4'b0000;
	ROM[2005] = 4'b0100;
	ROM[2006] = 4'b0000;
	ROM[2007] = 4'b1000;
	ROM[2008] = 4'b1100;
	ROM[2009] = 4'b1100;
	ROM[2010] = 4'b0000;
	ROM[2011] = 4'b0010;
	ROM[2012] = 4'b0011;
	ROM[2013] = 4'b0011;
	ROM[2014] = 4'b0000;
	ROM[2015] = 4'b0100;
	ROM[2016] = 4'b0000;
	ROM[2017] = 4'b0100;
	ROM[2018] = 4'b0000;
	ROM[2019] = 4'b0100;
	ROM[2020] = 4'b0000;
	ROM[2021] = 4'b0001;
	ROM[2022] = 4'b0000;
	ROM[2023] = 4'b0001;
	ROM[2024] = 4'b0000;
	ROM[2025] = 4'b0100;
	ROM[2026] = 4'b0000;
	ROM[2027] = 4'b0100;
	ROM[2028] = 4'b0000;
	ROM[2029] = 4'b0001;
	ROM[2030] = 4'b0000;
	ROM[2031] = 4'b0001;
	ROM[2032] = 4'b0000;
	ROM[2033] = 4'b0100;
	ROM[2034] = 4'b0000;
	ROM[2035] = 4'b0100;
	ROM[2036] = 4'b0000;
	ROM[2037] = 4'b0001;
	ROM[2038] = 4'b0000;
	ROM[2039] = 4'b0001;
	ROM[2040] = 4'b0000;
	ROM[2041] = 4'b0000;
	ROM[2042] = 4'b0000;
	ROM[2043] = 4'b0100;
	ROM[2044] = 4'b0000;
	ROM[2045] = 4'b0000;
	ROM[2046] = 4'b0000;
	ROM[2047] = 4'b0100;
	ROM[2048] = 4'b0000;
	ROM[2049] = 4'b1000;
	ROM[2050] = 4'b1100;
	ROM[2051] = 4'b1100;
	ROM[2052] = 4'b0000;
	ROM[2053] = 4'b0001;
	ROM[2054] = 4'b0000;
	ROM[2055] = 4'b0001;
	ROM[2056] = 4'b0000;
	ROM[2057] = 4'b0100;
	ROM[2058] = 4'b0000;
	ROM[2059] = 4'b0100;
	ROM[2060] = 4'b0000;
	ROM[2061] = 4'b0001;
	ROM[2062] = 4'b0000;
	ROM[2063] = 4'b0010;
	ROM[2064] = 4'b0011;
	ROM[2065] = 4'b0011;
	ROM[2066] = 4'b0000;
	ROM[2067] = 4'b0100;
	ROM[2068] = 4'b0000;
	ROM[2069] = 4'b0100;
	ROM[2070] = 4'b0000;
	ROM[2071] = 4'b1000;
	ROM[2072] = 4'b1100;
	ROM[2073] = 4'b1100;
	ROM[2074] = 4'b0000;
	ROM[2075] = 4'b0010;
	ROM[2076] = 4'b0011;
	ROM[2077] = 4'b0011;
	ROM[2078] = 4'b0000;
	ROM[2079] = 4'b0100;
	ROM[2080] = 4'b0000;
	ROM[2081] = 4'b0100;
	ROM[2082] = 4'b0000;
	ROM[2083] = 4'b0100;
	ROM[2084] = 4'b0000;
	ROM[2085] = 4'b0001;
	ROM[2086] = 4'b0000;
	ROM[2087] = 4'b0001;
	ROM[2088] = 4'b0000;
	ROM[2089] = 4'b0100;
	ROM[2090] = 4'b0000;
	ROM[2091] = 4'b0100;
	ROM[2092] = 4'b0000;
	ROM[2093] = 4'b0100;
	ROM[2094] = 4'b0000;
	ROM[2095] = 4'b0100;
	ROM[2096] = 4'b0000;
	ROM[2097] = 4'b0101;
	ROM[2098] = 4'b0000;
	ROM[2099] = 4'b0000;
	ROM[2100] = 4'b0000;
	ROM[2101] = 4'b0000;
	ROM[2102] = 4'b0000;
	ROM[2103] = 4'b0101;
	ROM[2104] = 4'b0000;
	ROM[2105] = 4'b0000;
	ROM[2106] = 4'b0000;
	ROM[2107] = 4'b0000;
	ROM[2108] = 4'b0000;
	ROM[2109] = 4'b0101;
	ROM[2110] = 4'b0000;
	ROM[2111] = 4'b0000;
	ROM[2112] = 4'b0000;
	ROM[2113] = 4'b0001;
	ROM[2114] = 4'b0000;
	ROM[2115] = 4'b0001;
	ROM[2116] = 4'b0000;
	ROM[2117] = 4'b0001;
	ROM[2118] = 4'b0000;
	ROM[2119] = 4'b0001;
	ROM[2120] = 4'b0000;
	ROM[2121] = 4'b0100;
	ROM[2122] = 4'b0000;
	ROM[2123] = 4'b0100;
	ROM[2124] = 4'b0000;
	ROM[2125] = 4'b0100;
	ROM[2126] = 4'b0000;
	ROM[2127] = 4'b0100;
	ROM[2128] = 4'b0000;
	ROM[2129] = 4'b0001;
	ROM[2130] = 4'b0000;
	ROM[2131] = 4'b0000;
	ROM[2132] = 4'b0001;
	ROM[2133] = 4'b0000;
	ROM[2134] = 4'b0000;
	ROM[2135] = 4'b0001;
	ROM[2136] = 4'b0000;
	ROM[2137] = 4'b0010;
	ROM[2138] = 4'b0011;
	ROM[2139] = 4'b0011;
	ROM[2140] = 4'b0011;
	ROM[2141] = 4'b0011;
	ROM[2142] = 4'b0000;
	ROM[2143] = 4'b0000;
	ROM[2144] = 4'b0000;
	ROM[2145] = 4'b0100;
	ROM[2146] = 4'b0000;
	ROM[2147] = 4'b0100;
	ROM[2148] = 4'b0000;
	ROM[2149] = 4'b0100;
	ROM[2150] = 4'b0000;
	ROM[2151] = 4'b0100;
	ROM[2152] = 4'b0000;
	ROM[2153] = 4'b0001;
	ROM[2154] = 4'b0000;
	ROM[2155] = 4'b0001;
	ROM[2156] = 4'b0000;
	ROM[2157] = 4'b0001;
	ROM[2158] = 4'b0000;
	ROM[2159] = 4'b0001;
	ROM[2160] = 4'b0000;
	ROM[2161] = 4'b0100;
	ROM[2162] = 4'b0000;
	ROM[2163] = 4'b0000;
	ROM[2164] = 4'b0100;
	ROM[2165] = 4'b0000;
	ROM[2166] = 4'b0000;
	ROM[2167] = 4'b0100;
	ROM[2168] = 4'b0000;
	ROM[2169] = 4'b1000;
	ROM[2170] = 4'b1100;
	ROM[2171] = 4'b1100;
	ROM[2172] = 4'b1100;
	ROM[2173] = 4'b1100;
	ROM[2174] = 4'b0000;
	ROM[2175] = 4'b0000;
	ROM[2176] = 4'b0000;
	ROM[2177] = 4'b0001;
	ROM[2178] = 4'b0000;
	ROM[2179] = 4'b0001;
	ROM[2180] = 4'b0000;
	ROM[2181] = 4'b0001;
	ROM[2182] = 4'b0000;
	ROM[2183] = 4'b0001;
	ROM[2184] = 4'b0000;
	ROM[2185] = 4'b0100;
	ROM[2186] = 4'b0000;
	ROM[2187] = 4'b0100;
	ROM[2188] = 4'b0000;
	ROM[2189] = 4'b0100;
	ROM[2190] = 4'b0000;
	ROM[2191] = 4'b0100;
	ROM[2192] = 4'b0000;
	ROM[2193] = 4'b0010;
	ROM[2194] = 4'b0011;
	ROM[2195] = 4'b0011;
	ROM[2196] = 4'b0011;
	ROM[2197] = 4'b0011;
	ROM[2198] = 4'b0011;
	ROM[2199] = 4'b0011;
	ROM[2200] = 4'b0011;
	ROM[2201] = 4'b1011;
	ROM[2202] = 4'b1100;
	ROM[2203] = 4'b1100;
	ROM[2204] = 4'b1100;
	ROM[2205] = 4'b1100;
	ROM[2206] = 4'b1100;
	ROM[2207] = 4'b1100;
	ROM[2208] = 4'b1100;
	ROM[2209] = 4'b1101;
	ROM[2210] = 4'b0000;
	ROM[2211] = 4'b0000;
	ROM[2212] = 4'b0000;
	ROM[2213] = 4'b0100;
	ROM[2214] = 4'b0000;
	ROM[2215] = 4'b0000;
	ROM[2216] = 4'b0000;
	ROM[2217] = 4'b0001;
	ROM[2218] = 4'b0000;
	ROM[2219] = 4'b0000;
	ROM[2220] = 4'b0000;
	ROM[2221] = 4'b0100;
	ROM[2222] = 4'b0000;
	ROM[2223] = 4'b0000;
	ROM[2224] = 4'b0000;
	ROM[2225] = 4'b1010;
	ROM[2226] = 4'b1111;
	ROM[2227] = 4'b1111;
	ROM[2228] = 4'b1111;
	ROM[2229] = 4'b1111;
	ROM[2230] = 4'b1111;
	ROM[2231] = 4'b1111;
	ROM[2232] = 4'b1111;
	ROM[2233] = 4'b1111;
	ROM[2234] = 4'b1111;
	ROM[2235] = 4'b1111;
	ROM[2236] = 4'b1111;
	ROM[2237] = 4'b1111;
	ROM[2238] = 4'b0000;
	ROM[2239] = 4'b0000;
	ROM[2240] = 4'b0000;
	ROM[2241] = 4'b0101;
	ROM[2242] = 4'b0000;
	ROM[2243] = 4'b0000;
	ROM[2244] = 4'b0000;
	ROM[2245] = 4'b0000;
	ROM[2246] = 4'b0000;
	ROM[2247] = 4'b0000;
	ROM[2248] = 4'b0000;
	ROM[2249] = 4'b0000;
	ROM[2250] = 4'b0000;
	ROM[2251] = 4'b0000;
	ROM[2252] = 4'b0000;
	ROM[2253] = 4'b0000;
	ROM[2254] = 4'b0000;
	ROM[2255] = 4'b0000;
	ROM[2256] = 4'b0000;
	ROM[2257] = 4'b0000;
	ROM[2258] = 4'b0000;
	ROM[2259] = 4'b0000;
	ROM[2260] = 4'b0000;
	ROM[2261] = 4'b0000;
	ROM[2262] = 4'b0000;
	ROM[2263] = 4'b0000;
	ROM[2264] = 4'b0000;
	ROM[2265] = 4'b0000;
	ROM[2266] = 4'b0000;
	ROM[2267] = 4'b0000;
	ROM[2268] = 4'b0000;
	ROM[2269] = 4'b0000;
	ROM[2270] = 4'b0000;
	ROM[2271] = 4'b0000;
	ROM[2272] = 4'b0000;
	ROM[2273] = 4'b0000;
	ROM[2274] = 4'b0000;
	ROM[2275] = 4'b0000;
	ROM[2276] = 4'b0000;
	ROM[2277] = 4'b0000;
	ROM[2278] = 4'b0000;
	ROM[2279] = 4'b0000;
	ROM[2280] = 4'b0000;
	ROM[2281] = 4'b0000;
	ROM[2282] = 4'b0000;
	ROM[2283] = 4'b0000;
	ROM[2284] = 4'b0000;
	ROM[2285] = 4'b0000;
	ROM[2286] = 4'b0000;
	ROM[2287] = 4'b0000;
	ROM[2288] = 4'b0000;
	ROM[2289] = 4'b0000;
	ROM[2290] = 4'b0000;
	ROM[2291] = 4'b0000;
	ROM[2292] = 4'b0000;
	ROM[2293] = 4'b0000;
	ROM[2294] = 4'b0000;
	ROM[2295] = 4'b0000;
	ROM[2296] = 4'b0000;
	ROM[2297] = 4'b0000;
	ROM[2298] = 4'b0000;
	ROM[2299] = 4'b0000;
	ROM[2300] = 4'b0000;
	ROM[2301] = 4'b0000;
	ROM[2302] = 4'b0000;
	ROM[2303] = 4'b0000;
	ROM[2304] = 4'b0000;
	ROM[2305] = 4'b0000;
	ROM[2306] = 4'b0000;
	ROM[2307] = 4'b0000;
	ROM[2308] = 4'b0000;
	ROM[2309] = 4'b0000;
	ROM[2310] = 4'b0000;
	ROM[2311] = 4'b0000;
	ROM[2312] = 4'b0000;
	ROM[2313] = 4'b0000;
	ROM[2314] = 4'b0000;
	ROM[2315] = 4'b0000;
	ROM[2316] = 4'b0000;
	ROM[2317] = 4'b0000;
	ROM[2318] = 4'b0000;
	ROM[2319] = 4'b0000;
	ROM[2320] = 4'b0000;
	ROM[2321] = 4'b0000;
	ROM[2322] = 4'b0000;
	ROM[2323] = 4'b0000;
	ROM[2324] = 4'b0000;
	ROM[2325] = 4'b0000;
	ROM[2326] = 4'b0000;
	ROM[2327] = 4'b0000;
	ROM[2328] = 4'b0000;
	ROM[2329] = 4'b0000;
	ROM[2330] = 4'b0000;
	ROM[2331] = 4'b0000;
	ROM[2332] = 4'b0000;
	ROM[2333] = 4'b0000;
	ROM[2334] = 4'b0000;
	ROM[2335] = 4'b0000;
	ROM[2336] = 4'b0000;
	ROM[2337] = 4'b0000;
	ROM[2338] = 4'b0000;
	ROM[2339] = 4'b0000;
	ROM[2340] = 4'b0000;
	ROM[2341] = 4'b0000;
	ROM[2342] = 4'b0000;
	ROM[2343] = 4'b0000;
	ROM[2344] = 4'b0000;
	ROM[2345] = 4'b0000;
	ROM[2346] = 4'b0000;
	ROM[2347] = 4'b0000;
	ROM[2348] = 4'b0000;
	ROM[2349] = 4'b0000;
	ROM[2350] = 4'b0000;
	ROM[2351] = 4'b0000;
	ROM[2352] = 4'b0000;
	ROM[2353] = 4'b0000;
	ROM[2354] = 4'b0000;
	ROM[2355] = 4'b0000;
	ROM[2356] = 4'b0000;
	ROM[2357] = 4'b0000;
	ROM[2358] = 4'b0000;
	ROM[2359] = 4'b0000;
	ROM[2360] = 4'b0000;
	ROM[2361] = 4'b0000;
	ROM[2362] = 4'b0000;
	ROM[2363] = 4'b0000;
	ROM[2364] = 4'b0000;
	ROM[2365] = 4'b0000;
	ROM[2366] = 4'b0000;
	ROM[2367] = 4'b0000;
	ROM[2368] = 4'b0000;
	ROM[2369] = 4'b0000;
	ROM[2370] = 4'b0000;
	ROM[2371] = 4'b0000;
	ROM[2372] = 4'b0000;
	ROM[2373] = 4'b0000;
	ROM[2374] = 4'b0000;
	ROM[2375] = 4'b0000;
	ROM[2376] = 4'b0000;
	ROM[2377] = 4'b0000;
	ROM[2378] = 4'b0000;
	ROM[2379] = 4'b0000;
	ROM[2380] = 4'b0000;
	ROM[2381] = 4'b0000;
	ROM[2382] = 4'b0000;
	ROM[2383] = 4'b0000;
	ROM[2384] = 4'b0000;
	ROM[2385] = 4'b0000;
	ROM[2386] = 4'b0000;
	ROM[2387] = 4'b0000;
	ROM[2388] = 4'b0000;
	ROM[2389] = 4'b0000;
	ROM[2390] = 4'b0000;
	ROM[2391] = 4'b0000;
	ROM[2392] = 4'b0000;
	ROM[2393] = 4'b0000;
	ROM[2394] = 4'b0000;
	ROM[2395] = 4'b0000;
	ROM[2396] = 4'b0000;
	ROM[2397] = 4'b0000;
	ROM[2398] = 4'b0000;
	ROM[2399] = 4'b0000;
	ROM[2400] = 4'b0000;
	ROM[2401] = 4'b0000;
	ROM[2402] = 4'b0000;
	ROM[2403] = 4'b0000;
	ROM[2404] = 4'b0000;
	ROM[2405] = 4'b0000;
	ROM[2406] = 4'b0000;
	ROM[2407] = 4'b0000;
	ROM[2408] = 4'b0000;
	ROM[2409] = 4'b0000;
	ROM[2410] = 4'b0000;
	ROM[2411] = 4'b0000;
	ROM[2412] = 4'b0000;
	ROM[2413] = 4'b0000;
	ROM[2414] = 4'b0000;
	ROM[2415] = 4'b0000;
	ROM[2416] = 4'b0000;
	ROM[2417] = 4'b0000;
	ROM[2418] = 4'b0000;
	ROM[2419] = 4'b0000;
	ROM[2420] = 4'b0000;
	ROM[2421] = 4'b0000;
	ROM[2422] = 4'b0000;
	ROM[2423] = 4'b0000;
	ROM[2424] = 4'b0000;
	ROM[2425] = 4'b0000;
	ROM[2426] = 4'b0000;
	ROM[2427] = 4'b0000;
	ROM[2428] = 4'b0000;
	ROM[2429] = 4'b0000;
	ROM[2430] = 4'b0000;
	ROM[2431] = 4'b0000;
	ROM[2432] = 4'b0000;
	ROM[2433] = 4'b0000;
	ROM[2434] = 4'b0000;
	ROM[2435] = 4'b0000;
	ROM[2436] = 4'b0000;
	ROM[2437] = 4'b0000;
	ROM[2438] = 4'b0000;
	ROM[2439] = 4'b0000;
	ROM[2440] = 4'b0000;
	ROM[2441] = 4'b0000;
	ROM[2442] = 4'b0000;
	ROM[2443] = 4'b0000;
	ROM[2444] = 4'b0000;
	ROM[2445] = 4'b0000;
	ROM[2446] = 4'b0000;
	ROM[2447] = 4'b0000;
	ROM[2448] = 4'b0000;
	ROM[2449] = 4'b0000;
	ROM[2450] = 4'b0000;
	ROM[2451] = 4'b0000;
	ROM[2452] = 4'b0000;
	ROM[2453] = 4'b0000;
	ROM[2454] = 4'b0000;
	ROM[2455] = 4'b0000;
	ROM[2456] = 4'b0000;
	ROM[2457] = 4'b0000;
	ROM[2458] = 4'b0000;
	ROM[2459] = 4'b0000;
	ROM[2460] = 4'b0000;
	ROM[2461] = 4'b0000;
	ROM[2462] = 4'b0000;
	ROM[2463] = 4'b0000;
	ROM[2464] = 4'b0000;
	ROM[2465] = 4'b0000;
	ROM[2466] = 4'b0000;
	ROM[2467] = 4'b0000;
	ROM[2468] = 4'b0000;
	ROM[2469] = 4'b0000;
	ROM[2470] = 4'b0000;
	ROM[2471] = 4'b0000;
	ROM[2472] = 4'b0000;
	ROM[2473] = 4'b0000;
	ROM[2474] = 4'b0000;
	ROM[2475] = 4'b0000;
	ROM[2476] = 4'b0000;
	ROM[2477] = 4'b0000;
	ROM[2478] = 4'b0000;
	ROM[2479] = 4'b0000;
	ROM[2480] = 4'b0000;
	ROM[2481] = 4'b0000;
	ROM[2482] = 4'b0000;
	ROM[2483] = 4'b0000;
	ROM[2484] = 4'b0000;
	ROM[2485] = 4'b0000;
	ROM[2486] = 4'b0000;
	ROM[2487] = 4'b0000;
	ROM[2488] = 4'b0000;
	ROM[2489] = 4'b0000;
	ROM[2490] = 4'b0000;
	ROM[2491] = 4'b0000;
	ROM[2492] = 4'b0000;
	ROM[2493] = 4'b0000;
	ROM[2494] = 4'b0000;
	ROM[2495] = 4'b0000;
	ROM[2496] = 4'b0000;
	ROM[2497] = 4'b0000;
	ROM[2498] = 4'b0000;
	ROM[2499] = 4'b0000;
	ROM[2500] = 4'b0000;
	ROM[2501] = 4'b0000;
	ROM[2502] = 4'b0000;
	ROM[2503] = 4'b0000;
	ROM[2504] = 4'b0000;
	ROM[2505] = 4'b0000;
	ROM[2506] = 4'b0000;
	ROM[2507] = 4'b0000;
	ROM[2508] = 4'b0000;
	ROM[2509] = 4'b0000;
	ROM[2510] = 4'b0000;
	ROM[2511] = 4'b0000;
	ROM[2512] = 4'b0000;
	ROM[2513] = 4'b0000;
	ROM[2514] = 4'b0000;
	ROM[2515] = 4'b0000;
	ROM[2516] = 4'b0000;
	ROM[2517] = 4'b0000;
	ROM[2518] = 4'b0000;
	ROM[2519] = 4'b0000;
	ROM[2520] = 4'b0000;
	ROM[2521] = 4'b0000;
	ROM[2522] = 4'b0000;
	ROM[2523] = 4'b0000;
	ROM[2524] = 4'b0000;
	ROM[2525] = 4'b0000;
	ROM[2526] = 4'b0000;
	ROM[2527] = 4'b0000;
	ROM[2528] = 4'b0000;
	ROM[2529] = 4'b0000;
	ROM[2530] = 4'b0000;
	ROM[2531] = 4'b0000;
	ROM[2532] = 4'b0000;
	ROM[2533] = 4'b0000;
	ROM[2534] = 4'b0000;
	ROM[2535] = 4'b0000;
	ROM[2536] = 4'b0000;
	ROM[2537] = 4'b0000;
	ROM[2538] = 4'b0000;
	ROM[2539] = 4'b0000;
	ROM[2540] = 4'b0000;
	ROM[2541] = 4'b0000;
	ROM[2542] = 4'b0000;
	ROM[2543] = 4'b0000;
	ROM[2544] = 4'b0000;
	ROM[2545] = 4'b0000;
	ROM[2546] = 4'b0000;
	ROM[2547] = 4'b0000;
	ROM[2548] = 4'b0000;
	ROM[2549] = 4'b0000;
	ROM[2550] = 4'b0000;
	ROM[2551] = 4'b0000;
	ROM[2552] = 4'b0000;
	ROM[2553] = 4'b0000;
	ROM[2554] = 4'b0000;
	ROM[2555] = 4'b0000;
	ROM[2556] = 4'b0000;
	ROM[2557] = 4'b0000;
	ROM[2558] = 4'b0000;
	ROM[2559] = 4'b0000;
	ROM[2560] = 4'b0000;
	ROM[2561] = 4'b0000;
	ROM[2562] = 4'b0000;
	ROM[2563] = 4'b0000;
	ROM[2564] = 4'b0000;
	ROM[2565] = 4'b0000;
	ROM[2566] = 4'b0000;
	ROM[2567] = 4'b0000;
	ROM[2568] = 4'b0000;
	ROM[2569] = 4'b0000;
	ROM[2570] = 4'b0000;
	ROM[2571] = 4'b0000;
	ROM[2572] = 4'b0000;
	ROM[2573] = 4'b0000;
	ROM[2574] = 4'b0000;
	ROM[2575] = 4'b0000;
	ROM[2576] = 4'b0000;
	ROM[2577] = 4'b0000;
	ROM[2578] = 4'b0000;
	ROM[2579] = 4'b0000;
	ROM[2580] = 4'b0000;
	ROM[2581] = 4'b0000;
	ROM[2582] = 4'b0000;
	ROM[2583] = 4'b0000;
	ROM[2584] = 4'b0000;
	ROM[2585] = 4'b0000;
	ROM[2586] = 4'b0000;
	ROM[2587] = 4'b0000;
	ROM[2588] = 4'b0000;
	ROM[2589] = 4'b0000;
	ROM[2590] = 4'b0000;
	ROM[2591] = 4'b0000;
	ROM[2592] = 4'b0000;
	ROM[2593] = 4'b0000;
	ROM[2594] = 4'b0000;
	ROM[2595] = 4'b0000;
	ROM[2596] = 4'b0000;
	ROM[2597] = 4'b0000;
	ROM[2598] = 4'b0000;
	ROM[2599] = 4'b0000;
	ROM[2600] = 4'b0000;
	ROM[2601] = 4'b0000;
	ROM[2602] = 4'b0000;
	ROM[2603] = 4'b0000;
	ROM[2604] = 4'b0000;
	ROM[2605] = 4'b0000;
	ROM[2606] = 4'b0000;
	ROM[2607] = 4'b0000;
	ROM[2608] = 4'b0000;
	ROM[2609] = 4'b0000;
	ROM[2610] = 4'b0000;
	ROM[2611] = 4'b0000;
	ROM[2612] = 4'b0000;
	ROM[2613] = 4'b0000;
	ROM[2614] = 4'b0000;
	ROM[2615] = 4'b0000;
	ROM[2616] = 4'b0000;
	ROM[2617] = 4'b0000;
	ROM[2618] = 4'b0000;
	ROM[2619] = 4'b0000;
	ROM[2620] = 4'b0000;
	ROM[2621] = 4'b0000;
	ROM[2622] = 4'b0000;
	ROM[2623] = 4'b0000;
	ROM[2624] = 4'b0000;
	ROM[2625] = 4'b0000;
	ROM[2626] = 4'b0000;
	ROM[2627] = 4'b0000;
	ROM[2628] = 4'b0000;
	ROM[2629] = 4'b0000;
	ROM[2630] = 4'b0000;
	ROM[2631] = 4'b0000;
	ROM[2632] = 4'b0000;
	ROM[2633] = 4'b0000;
	ROM[2634] = 4'b0000;
	ROM[2635] = 4'b0000;
	ROM[2636] = 4'b0000;
	ROM[2637] = 4'b0000;
	ROM[2638] = 4'b0000;
	ROM[2639] = 4'b0000;
	ROM[2640] = 4'b0000;
	ROM[2641] = 4'b0000;
	ROM[2642] = 4'b0000;
	ROM[2643] = 4'b0000;
	ROM[2644] = 4'b0000;
	ROM[2645] = 4'b0000;
	ROM[2646] = 4'b0000;
	ROM[2647] = 4'b0000;
	ROM[2648] = 4'b0000;
	ROM[2649] = 4'b0000;
	ROM[2650] = 4'b0000;
	ROM[2651] = 4'b0000;
	ROM[2652] = 4'b0000;
	ROM[2653] = 4'b0000;
	ROM[2654] = 4'b0000;
	ROM[2655] = 4'b0000;
	ROM[2656] = 4'b0000;
	ROM[2657] = 4'b0000;
	ROM[2658] = 4'b0000;
	ROM[2659] = 4'b0000;
	ROM[2660] = 4'b0000;
	ROM[2661] = 4'b0000;
	ROM[2662] = 4'b0000;
	ROM[2663] = 4'b0000;
	ROM[2664] = 4'b0000;
	ROM[2665] = 4'b0000;
	ROM[2666] = 4'b0000;
	ROM[2667] = 4'b0000;
	ROM[2668] = 4'b0000;
	ROM[2669] = 4'b0000;
	ROM[2670] = 4'b0000;
	ROM[2671] = 4'b0000;
	ROM[2672] = 4'b0000;
	ROM[2673] = 4'b0000;
	ROM[2674] = 4'b0000;
	ROM[2675] = 4'b0000;
	ROM[2676] = 4'b0000;
	ROM[2677] = 4'b0000;
	ROM[2678] = 4'b0000;
	ROM[2679] = 4'b0000;
	ROM[2680] = 4'b0000;
	ROM[2681] = 4'b0000;
	ROM[2682] = 4'b0000;
	ROM[2683] = 4'b0000;
	ROM[2684] = 4'b0000;
	ROM[2685] = 4'b0000;
	ROM[2686] = 4'b0000;
	ROM[2687] = 4'b0000;
	ROM[2688] = 4'b0000;
	ROM[2689] = 4'b0000;
	ROM[2690] = 4'b0000;
	ROM[2691] = 4'b0000;
	ROM[2692] = 4'b0000;
	ROM[2693] = 4'b0000;
	ROM[2694] = 4'b0000;
	ROM[2695] = 4'b0000;
	ROM[2696] = 4'b0000;
	ROM[2697] = 4'b0000;
	ROM[2698] = 4'b0000;
	ROM[2699] = 4'b0000;
	ROM[2700] = 4'b0000;
	ROM[2701] = 4'b0000;
	ROM[2702] = 4'b0000;
	ROM[2703] = 4'b0000;
	ROM[2704] = 4'b0000;
	ROM[2705] = 4'b0000;
	ROM[2706] = 4'b0000;
	ROM[2707] = 4'b0000;
	ROM[2708] = 4'b0000;
	ROM[2709] = 4'b0000;
	ROM[2710] = 4'b0000;
	ROM[2711] = 4'b0000;
	ROM[2712] = 4'b0000;
	ROM[2713] = 4'b0000;
	ROM[2714] = 4'b0000;
	ROM[2715] = 4'b0000;
	ROM[2716] = 4'b0000;
	ROM[2717] = 4'b0000;
	ROM[2718] = 4'b0000;
	ROM[2719] = 4'b0000;
	ROM[2720] = 4'b0000;
	ROM[2721] = 4'b0000;
	ROM[2722] = 4'b0000;
	ROM[2723] = 4'b0000;
	ROM[2724] = 4'b0000;
	ROM[2725] = 4'b0000;
	ROM[2726] = 4'b0000;
	ROM[2727] = 4'b0000;
	ROM[2728] = 4'b0000;
	ROM[2729] = 4'b0000;
	ROM[2730] = 4'b0000;
	ROM[2731] = 4'b0000;
	ROM[2732] = 4'b0000;
	ROM[2733] = 4'b0000;
	ROM[2734] = 4'b0000;
	ROM[2735] = 4'b0000;
	ROM[2736] = 4'b0000;
	ROM[2737] = 4'b0000;
	ROM[2738] = 4'b0000;
	ROM[2739] = 4'b0000;
	ROM[2740] = 4'b0000;
	ROM[2741] = 4'b0000;
	ROM[2742] = 4'b0000;
	ROM[2743] = 4'b0000;
	ROM[2744] = 4'b0000;
	ROM[2745] = 4'b0000;
	ROM[2746] = 4'b0000;
	ROM[2747] = 4'b0000;
	ROM[2748] = 4'b0000;
	ROM[2749] = 4'b0000;
	ROM[2750] = 4'b0000;
	ROM[2751] = 4'b0000;
	ROM[2752] = 4'b0000;
	ROM[2753] = 4'b0000;
	ROM[2754] = 4'b0000;
	ROM[2755] = 4'b0000;
	ROM[2756] = 4'b0000;
	ROM[2757] = 4'b0000;
	ROM[2758] = 4'b0000;
	ROM[2759] = 4'b0000;
	ROM[2760] = 4'b0000;
	ROM[2761] = 4'b0000;
	ROM[2762] = 4'b0000;
	ROM[2763] = 4'b0000;
	ROM[2764] = 4'b0000;
	ROM[2765] = 4'b0000;
	ROM[2766] = 4'b0000;
	ROM[2767] = 4'b0000;
	ROM[2768] = 4'b0000;
	ROM[2769] = 4'b0000;
	ROM[2770] = 4'b0000;
	ROM[2771] = 4'b0000;
	ROM[2772] = 4'b0000;
	ROM[2773] = 4'b0000;
	ROM[2774] = 4'b0000;
	ROM[2775] = 4'b0000;
	ROM[2776] = 4'b0000;
	ROM[2777] = 4'b0000;
	ROM[2778] = 4'b0000;
	ROM[2779] = 4'b0000;
	ROM[2780] = 4'b0000;
	ROM[2781] = 4'b0000;
	ROM[2782] = 4'b0000;
	ROM[2783] = 4'b0000;
	ROM[2784] = 4'b0000;
	ROM[2785] = 4'b0000;
	ROM[2786] = 4'b0000;
	ROM[2787] = 4'b0000;
	ROM[2788] = 4'b0000;
	ROM[2789] = 4'b0000;
	ROM[2790] = 4'b0000;
	ROM[2791] = 4'b0000;
	ROM[2792] = 4'b0000;
	ROM[2793] = 4'b0000;
	ROM[2794] = 4'b0000;
	ROM[2795] = 4'b0000;
	ROM[2796] = 4'b0000;
	ROM[2797] = 4'b0000;
	ROM[2798] = 4'b0000;
	ROM[2799] = 4'b0000;
	ROM[2800] = 4'b0000;
	ROM[2801] = 4'b0000;
	ROM[2802] = 4'b0000;
	ROM[2803] = 4'b0000;
	ROM[2804] = 4'b0000;
	ROM[2805] = 4'b0000;
	ROM[2806] = 4'b0000;
	ROM[2807] = 4'b0000;
	ROM[2808] = 4'b0000;
	ROM[2809] = 4'b0000;
	ROM[2810] = 4'b0000;
	ROM[2811] = 4'b0000;
	ROM[2812] = 4'b0000;
	ROM[2813] = 4'b0000;
	ROM[2814] = 4'b0000;
	ROM[2815] = 4'b0000;
	ROM[2816] = 4'b0000;
	ROM[2817] = 4'b0000;
	ROM[2818] = 4'b0000;
	ROM[2819] = 4'b0000;
	ROM[2820] = 4'b0000;
	ROM[2821] = 4'b0000;
	ROM[2822] = 4'b0000;
	ROM[2823] = 4'b0000;
	ROM[2824] = 4'b0000;
	ROM[2825] = 4'b0000;
	ROM[2826] = 4'b0000;
	ROM[2827] = 4'b0000;
	ROM[2828] = 4'b0000;
	ROM[2829] = 4'b0000;
	ROM[2830] = 4'b0000;
	ROM[2831] = 4'b0000;
	ROM[2832] = 4'b0000;
	ROM[2833] = 4'b0000;
	ROM[2834] = 4'b0000;
	ROM[2835] = 4'b0000;
	ROM[2836] = 4'b0000;
	ROM[2837] = 4'b0000;
	ROM[2838] = 4'b0000;
	ROM[2839] = 4'b0000;
	ROM[2840] = 4'b0000;
	ROM[2841] = 4'b0000;
	ROM[2842] = 4'b0000;
	ROM[2843] = 4'b0000;
	ROM[2844] = 4'b0000;
	ROM[2845] = 4'b0000;
	ROM[2846] = 4'b0000;
	ROM[2847] = 4'b0000;
	ROM[2848] = 4'b0000;
	ROM[2849] = 4'b0000;
	ROM[2850] = 4'b0000;
	ROM[2851] = 4'b0000;
	ROM[2852] = 4'b0000;
	ROM[2853] = 4'b0000;
	ROM[2854] = 4'b0000;
	ROM[2855] = 4'b0000;
	ROM[2856] = 4'b0000;
	ROM[2857] = 4'b0000;
	ROM[2858] = 4'b0000;
	ROM[2859] = 4'b0000;
	ROM[2860] = 4'b0000;
	ROM[2861] = 4'b0000;
	ROM[2862] = 4'b0000;
	ROM[2863] = 4'b0000;
	ROM[2864] = 4'b0000;
	ROM[2865] = 4'b0000;
	ROM[2866] = 4'b0000;
	ROM[2867] = 4'b0000;
	ROM[2868] = 4'b0000;
	ROM[2869] = 4'b0000;
	ROM[2870] = 4'b0000;
	ROM[2871] = 4'b0000;
	ROM[2872] = 4'b0000;
	ROM[2873] = 4'b0000;
	ROM[2874] = 4'b0000;
	ROM[2875] = 4'b0000;
	ROM[2876] = 4'b0000;
	ROM[2877] = 4'b0000;
	ROM[2878] = 4'b0000;
	ROM[2879] = 4'b0000;
	ROM[2880] = 4'b0000;
	ROM[2881] = 4'b0000;
	ROM[2882] = 4'b0000;
	ROM[2883] = 4'b0000;
	ROM[2884] = 4'b0000;
	ROM[2885] = 4'b0000;
	ROM[2886] = 4'b0000;
	ROM[2887] = 4'b0000;
	ROM[2888] = 4'b0000;
	ROM[2889] = 4'b0000;
	ROM[2890] = 4'b0000;
	ROM[2891] = 4'b0000;
	ROM[2892] = 4'b0000;
	ROM[2893] = 4'b0000;
	ROM[2894] = 4'b0000;
	ROM[2895] = 4'b0000;
	ROM[2896] = 4'b0000;
	ROM[2897] = 4'b0000;
	ROM[2898] = 4'b0000;
	ROM[2899] = 4'b0000;
	ROM[2900] = 4'b0000;
	ROM[2901] = 4'b0000;
	ROM[2902] = 4'b0000;
	ROM[2903] = 4'b0000;
	ROM[2904] = 4'b0000;
	ROM[2905] = 4'b0000;
	ROM[2906] = 4'b0000;
	ROM[2907] = 4'b0000;
	ROM[2908] = 4'b0000;
	ROM[2909] = 4'b0000;
	ROM[2910] = 4'b0000;
	ROM[2911] = 4'b0000;
	ROM[2912] = 4'b0000;
	ROM[2913] = 4'b0000;
	ROM[2914] = 4'b0000;
	ROM[2915] = 4'b0000;
	ROM[2916] = 4'b0000;
	ROM[2917] = 4'b0000;
	ROM[2918] = 4'b0000;
	ROM[2919] = 4'b0000;
	ROM[2920] = 4'b0000;
	ROM[2921] = 4'b0000;
	ROM[2922] = 4'b0000;
	ROM[2923] = 4'b0000;
	ROM[2924] = 4'b0000;
	ROM[2925] = 4'b0000;
	ROM[2926] = 4'b0000;
	ROM[2927] = 4'b0000;
	ROM[2928] = 4'b0000;
	ROM[2929] = 4'b0000;
	ROM[2930] = 4'b0000;
	ROM[2931] = 4'b0000;
	ROM[2932] = 4'b0000;
	ROM[2933] = 4'b0000;
	ROM[2934] = 4'b0000;
	ROM[2935] = 4'b0000;
	ROM[2936] = 4'b0000;
	ROM[2937] = 4'b0000;
	ROM[2938] = 4'b0000;
	ROM[2939] = 4'b0000;
	ROM[2940] = 4'b0000;
	ROM[2941] = 4'b0000;
	ROM[2942] = 4'b0000;
	ROM[2943] = 4'b0000;
	ROM[2944] = 4'b0000;
	ROM[2945] = 4'b0000;
	ROM[2946] = 4'b0000;
	ROM[2947] = 4'b0000;
	ROM[2948] = 4'b0000;
	ROM[2949] = 4'b0000;
	ROM[2950] = 4'b0000;
	ROM[2951] = 4'b0000;
	ROM[2952] = 4'b0000;
	ROM[2953] = 4'b0000;
	ROM[2954] = 4'b0000;
	ROM[2955] = 4'b0000;
	ROM[2956] = 4'b0000;
	ROM[2957] = 4'b0000;
	ROM[2958] = 4'b0000;
	ROM[2959] = 4'b0000;
	ROM[2960] = 4'b0000;
	ROM[2961] = 4'b0000;
	ROM[2962] = 4'b0000;
	ROM[2963] = 4'b0000;
	ROM[2964] = 4'b0000;
	ROM[2965] = 4'b0000;
	ROM[2966] = 4'b0000;
	ROM[2967] = 4'b0000;
	ROM[2968] = 4'b0000;
	ROM[2969] = 4'b0000;
	ROM[2970] = 4'b0000;
	ROM[2971] = 4'b0000;
	ROM[2972] = 4'b0000;
	ROM[2973] = 4'b0000;
	ROM[2974] = 4'b0000;
	ROM[2975] = 4'b0000;
	ROM[2976] = 4'b0000;
	ROM[2977] = 4'b0000;
	ROM[2978] = 4'b0000;
	ROM[2979] = 4'b0000;
	ROM[2980] = 4'b0000;
	ROM[2981] = 4'b0000;
	ROM[2982] = 4'b0000;
	ROM[2983] = 4'b0000;
	ROM[2984] = 4'b0000;
	ROM[2985] = 4'b0000;
	ROM[2986] = 4'b0000;
	ROM[2987] = 4'b0000;
	ROM[2988] = 4'b0000;
	ROM[2989] = 4'b0000;
	ROM[2990] = 4'b0000;
	ROM[2991] = 4'b0000;
	ROM[2992] = 4'b0000;
	ROM[2993] = 4'b0000;
	ROM[2994] = 4'b0000;
	ROM[2995] = 4'b0000;
	ROM[2996] = 4'b0000;
	ROM[2997] = 4'b0000;
	ROM[2998] = 4'b0000;
	ROM[2999] = 4'b0000;
	ROM[3000] = 4'b0000;
	ROM[3001] = 4'b0000;
	ROM[3002] = 4'b0000;
	ROM[3003] = 4'b0000;
	ROM[3004] = 4'b0000;
	ROM[3005] = 4'b0000;
	ROM[3006] = 4'b0000;
	ROM[3007] = 4'b0000;
	ROM[3008] = 4'b0000;
	ROM[3009] = 4'b0000;
	ROM[3010] = 4'b0000;
	ROM[3011] = 4'b0000;
	ROM[3012] = 4'b0000;
	ROM[3013] = 4'b0000;
	ROM[3014] = 4'b0000;
	ROM[3015] = 4'b0000;
	ROM[3016] = 4'b0000;
	ROM[3017] = 4'b0000;
	ROM[3018] = 4'b0000;
	ROM[3019] = 4'b0000;
	ROM[3020] = 4'b0000;
	ROM[3021] = 4'b0000;
	ROM[3022] = 4'b0000;
	ROM[3023] = 4'b0000;
	ROM[3024] = 4'b0000;
	ROM[3025] = 4'b0000;
	ROM[3026] = 4'b0000;
	ROM[3027] = 4'b0000;
	ROM[3028] = 4'b0000;
	ROM[3029] = 4'b0000;
	ROM[3030] = 4'b0000;
	ROM[3031] = 4'b0000;
	ROM[3032] = 4'b0000;
	ROM[3033] = 4'b0000;
	ROM[3034] = 4'b0000;
	ROM[3035] = 4'b0000;
	ROM[3036] = 4'b0000;
	ROM[3037] = 4'b0000;
	ROM[3038] = 4'b0000;
	ROM[3039] = 4'b0000;
	ROM[3040] = 4'b0000;
	ROM[3041] = 4'b0000;
	ROM[3042] = 4'b0000;
	ROM[3043] = 4'b0000;
	ROM[3044] = 4'b0000;
	ROM[3045] = 4'b0000;
	ROM[3046] = 4'b0000;
	ROM[3047] = 4'b0000;
	ROM[3048] = 4'b0000;
	ROM[3049] = 4'b0000;
	ROM[3050] = 4'b0000;
	ROM[3051] = 4'b0000;
	ROM[3052] = 4'b0000;
	ROM[3053] = 4'b0000;
	ROM[3054] = 4'b0000;
	ROM[3055] = 4'b0000;
	ROM[3056] = 4'b0000;
	ROM[3057] = 4'b0000;
	ROM[3058] = 4'b0000;
	ROM[3059] = 4'b0000;
	ROM[3060] = 4'b0000;
	ROM[3061] = 4'b0000;
	ROM[3062] = 4'b0000;
	ROM[3063] = 4'b0000;
	ROM[3064] = 4'b0000;
	ROM[3065] = 4'b0000;
	ROM[3066] = 4'b0000;
	ROM[3067] = 4'b0000;
	ROM[3068] = 4'b0000;
	ROM[3069] = 4'b0000;
	ROM[3070] = 4'b0000;
	ROM[3071] = 4'b0000;
	ROM[3072] = 4'b0000;
	ROM[3073] = 4'b0000;
	ROM[3074] = 4'b0000;
	ROM[3075] = 4'b0000;
	ROM[3076] = 4'b0000;
	ROM[3077] = 4'b0000;
	ROM[3078] = 4'b0000;
	ROM[3079] = 4'b0000;
	ROM[3080] = 4'b0000;
	ROM[3081] = 4'b0000;
	ROM[3082] = 4'b0000;
	ROM[3083] = 4'b0000;
	ROM[3084] = 4'b0000;
	ROM[3085] = 4'b0000;
	ROM[3086] = 4'b0000;
	ROM[3087] = 4'b0000;
	ROM[3088] = 4'b0000;
	ROM[3089] = 4'b0000;
	ROM[3090] = 4'b0000;
	ROM[3091] = 4'b0000;
	ROM[3092] = 4'b0000;
	ROM[3093] = 4'b0000;
	ROM[3094] = 4'b0000;
	ROM[3095] = 4'b0000;
	ROM[3096] = 4'b0000;
	ROM[3097] = 4'b0000;
	ROM[3098] = 4'b0000;
	ROM[3099] = 4'b0000;
	ROM[3100] = 4'b0000;
	ROM[3101] = 4'b0000;
	ROM[3102] = 4'b0000;
	ROM[3103] = 4'b0000;
	ROM[3104] = 4'b0000;
	ROM[3105] = 4'b0000;
	ROM[3106] = 4'b0000;
	ROM[3107] = 4'b0000;
	ROM[3108] = 4'b0000;
	ROM[3109] = 4'b0000;
	ROM[3110] = 4'b0000;
	ROM[3111] = 4'b0000;
	ROM[3112] = 4'b0000;
	ROM[3113] = 4'b0000;
	ROM[3114] = 4'b0000;
	ROM[3115] = 4'b0000;
	ROM[3116] = 4'b0000;
	ROM[3117] = 4'b0000;
	ROM[3118] = 4'b0000;
	ROM[3119] = 4'b0000;
	ROM[3120] = 4'b0000;
	ROM[3121] = 4'b0000;
	ROM[3122] = 4'b0000;
	ROM[3123] = 4'b0000;
	ROM[3124] = 4'b0000;
	ROM[3125] = 4'b0000;
	ROM[3126] = 4'b0000;
	ROM[3127] = 4'b0000;
	ROM[3128] = 4'b0000;
	ROM[3129] = 4'b0000;
	ROM[3130] = 4'b0000;
	ROM[3131] = 4'b0000;
	ROM[3132] = 4'b0000;
	ROM[3133] = 4'b0000;
	ROM[3134] = 4'b0000;
	ROM[3135] = 4'b0000;
	ROM[3136] = 4'b0000;
	ROM[3137] = 4'b0000;
	ROM[3138] = 4'b0000;
	ROM[3139] = 4'b0000;
	ROM[3140] = 4'b0000;
	ROM[3141] = 4'b0000;
	ROM[3142] = 4'b0000;
	ROM[3143] = 4'b0000;
	ROM[3144] = 4'b0000;
	ROM[3145] = 4'b0000;
	ROM[3146] = 4'b0000;
	ROM[3147] = 4'b0000;
	ROM[3148] = 4'b0000;
	ROM[3149] = 4'b0000;
	ROM[3150] = 4'b0000;
	ROM[3151] = 4'b0000;
	ROM[3152] = 4'b0000;
	ROM[3153] = 4'b0000;
	ROM[3154] = 4'b0000;
	ROM[3155] = 4'b0000;
	ROM[3156] = 4'b0000;
	ROM[3157] = 4'b0000;
	ROM[3158] = 4'b0000;
	ROM[3159] = 4'b0000;
	ROM[3160] = 4'b0000;
	ROM[3161] = 4'b0000;
	ROM[3162] = 4'b0000;
	ROM[3163] = 4'b0000;
	ROM[3164] = 4'b0000;
	ROM[3165] = 4'b0000;
	ROM[3166] = 4'b0000;
	ROM[3167] = 4'b0000;
	ROM[3168] = 4'b0000;
	ROM[3169] = 4'b0000;
	ROM[3170] = 4'b0000;
	ROM[3171] = 4'b0000;
	ROM[3172] = 4'b0000;
	ROM[3173] = 4'b0000;
	ROM[3174] = 4'b0000;
	ROM[3175] = 4'b0000;
	ROM[3176] = 4'b0000;
	ROM[3177] = 4'b0000;
	ROM[3178] = 4'b0000;
	ROM[3179] = 4'b0000;
	ROM[3180] = 4'b0000;
	ROM[3181] = 4'b0000;
	ROM[3182] = 4'b0000;
	ROM[3183] = 4'b0000;
	ROM[3184] = 4'b0000;
	ROM[3185] = 4'b0000;
	ROM[3186] = 4'b0000;
	ROM[3187] = 4'b0000;
	ROM[3188] = 4'b0000;
	ROM[3189] = 4'b0000;
	ROM[3190] = 4'b0000;
	ROM[3191] = 4'b0000;
	ROM[3192] = 4'b0000;
	ROM[3193] = 4'b0000;
	ROM[3194] = 4'b0000;
	ROM[3195] = 4'b0000;
	ROM[3196] = 4'b0000;
	ROM[3197] = 4'b0000;
	ROM[3198] = 4'b0000;
	ROM[3199] = 4'b0000;
	ROM[3200] = 4'b0000;
	ROM[3201] = 4'b0000;
	ROM[3202] = 4'b0000;
	ROM[3203] = 4'b0000;
	ROM[3204] = 4'b0000;
	ROM[3205] = 4'b0000;
	ROM[3206] = 4'b0000;
	ROM[3207] = 4'b0000;
	ROM[3208] = 4'b0000;
	ROM[3209] = 4'b0000;
	ROM[3210] = 4'b0000;
	ROM[3211] = 4'b0000;
	ROM[3212] = 4'b0000;
	ROM[3213] = 4'b0000;
	ROM[3214] = 4'b0000;
	ROM[3215] = 4'b0000;
	ROM[3216] = 4'b0000;
	ROM[3217] = 4'b0000;
	ROM[3218] = 4'b0000;
	ROM[3219] = 4'b0000;
	ROM[3220] = 4'b0000;
	ROM[3221] = 4'b0000;
	ROM[3222] = 4'b0000;
	ROM[3223] = 4'b0000;
	ROM[3224] = 4'b0000;
	ROM[3225] = 4'b0000;
	ROM[3226] = 4'b0000;
	ROM[3227] = 4'b0000;
	ROM[3228] = 4'b0000;
	ROM[3229] = 4'b0000;
	ROM[3230] = 4'b0000;
	ROM[3231] = 4'b0000;
	ROM[3232] = 4'b0000;
	ROM[3233] = 4'b0000;
	ROM[3234] = 4'b0000;
	ROM[3235] = 4'b0000;
	ROM[3236] = 4'b0000;
	ROM[3237] = 4'b0000;
	ROM[3238] = 4'b0000;
	ROM[3239] = 4'b0000;
	ROM[3240] = 4'b0000;
	ROM[3241] = 4'b0000;
	ROM[3242] = 4'b0000;
	ROM[3243] = 4'b0000;
	ROM[3244] = 4'b0000;
	ROM[3245] = 4'b0000;
	ROM[3246] = 4'b0000;
	ROM[3247] = 4'b0000;
	ROM[3248] = 4'b0000;
	ROM[3249] = 4'b0000;
	ROM[3250] = 4'b0000;
	ROM[3251] = 4'b0000;
	ROM[3252] = 4'b0000;
	ROM[3253] = 4'b0000;
	ROM[3254] = 4'b0000;
	ROM[3255] = 4'b0000;
	ROM[3256] = 4'b0000;
	ROM[3257] = 4'b0000;
	ROM[3258] = 4'b0000;
	ROM[3259] = 4'b0000;
	ROM[3260] = 4'b0000;
	ROM[3261] = 4'b0000;
	ROM[3262] = 4'b0000;
	ROM[3263] = 4'b0000;
	ROM[3264] = 4'b0000;
	ROM[3265] = 4'b0000;
	ROM[3266] = 4'b0000;
	ROM[3267] = 4'b0000;
	ROM[3268] = 4'b0000;
	ROM[3269] = 4'b0000;
	ROM[3270] = 4'b0000;
	ROM[3271] = 4'b0000;
	ROM[3272] = 4'b0000;
	ROM[3273] = 4'b0000;
	ROM[3274] = 4'b0000;
	ROM[3275] = 4'b0000;
	ROM[3276] = 4'b0000;
	ROM[3277] = 4'b0000;
	ROM[3278] = 4'b0000;
	ROM[3279] = 4'b0000;
	ROM[3280] = 4'b0000;
	ROM[3281] = 4'b0000;
	ROM[3282] = 4'b0000;
	ROM[3283] = 4'b0000;
	ROM[3284] = 4'b0000;
	ROM[3285] = 4'b0000;
	ROM[3286] = 4'b0000;
	ROM[3287] = 4'b0000;
	ROM[3288] = 4'b0000;
	ROM[3289] = 4'b0000;
	ROM[3290] = 4'b0000;
	ROM[3291] = 4'b0000;
	ROM[3292] = 4'b0000;
	ROM[3293] = 4'b0000;
	ROM[3294] = 4'b0000;
	ROM[3295] = 4'b0000;
	ROM[3296] = 4'b0000;
	ROM[3297] = 4'b0000;
	ROM[3298] = 4'b0000;
	ROM[3299] = 4'b0000;
	ROM[3300] = 4'b0000;
	ROM[3301] = 4'b0000;
	ROM[3302] = 4'b0000;
	ROM[3303] = 4'b0000;
	ROM[3304] = 4'b0000;
	ROM[3305] = 4'b0000;
	ROM[3306] = 4'b0000;
	ROM[3307] = 4'b0000;
	ROM[3308] = 4'b0000;
	ROM[3309] = 4'b0000;
	ROM[3310] = 4'b0000;
	ROM[3311] = 4'b0000;
	ROM[3312] = 4'b0000;
	ROM[3313] = 4'b0000;
	ROM[3314] = 4'b0000;
	ROM[3315] = 4'b0000;
	ROM[3316] = 4'b0000;
	ROM[3317] = 4'b0000;
	ROM[3318] = 4'b0000;
	ROM[3319] = 4'b0000;
	ROM[3320] = 4'b0000;
	ROM[3321] = 4'b0000;
	ROM[3322] = 4'b0000;
	ROM[3323] = 4'b0000;
	ROM[3324] = 4'b0000;
	ROM[3325] = 4'b0000;
	ROM[3326] = 4'b0000;
	ROM[3327] = 4'b0000;
	ROM[3328] = 4'b0000;
	ROM[3329] = 4'b0000;
	ROM[3330] = 4'b0000;
	ROM[3331] = 4'b0000;
	ROM[3332] = 4'b0000;
	ROM[3333] = 4'b0000;
	ROM[3334] = 4'b0000;
	ROM[3335] = 4'b0000;
	ROM[3336] = 4'b0000;
	ROM[3337] = 4'b0000;
	ROM[3338] = 4'b0000;
	ROM[3339] = 4'b0000;
	ROM[3340] = 4'b0000;
	ROM[3341] = 4'b0000;
	ROM[3342] = 4'b0000;
	ROM[3343] = 4'b0000;
	ROM[3344] = 4'b0000;
	ROM[3345] = 4'b0000;
	ROM[3346] = 4'b0000;
	ROM[3347] = 4'b0000;
	ROM[3348] = 4'b0000;
	ROM[3349] = 4'b0000;
	ROM[3350] = 4'b0000;
	ROM[3351] = 4'b0000;
	ROM[3352] = 4'b0000;
	ROM[3353] = 4'b0000;
	ROM[3354] = 4'b0000;
	ROM[3355] = 4'b0000;
	ROM[3356] = 4'b0000;
	ROM[3357] = 4'b0000;
	ROM[3358] = 4'b0000;
	ROM[3359] = 4'b0000;
	ROM[3360] = 4'b0000;
	ROM[3361] = 4'b0000;
	ROM[3362] = 4'b0000;
	ROM[3363] = 4'b0000;
	ROM[3364] = 4'b0000;
	ROM[3365] = 4'b0000;
	ROM[3366] = 4'b0000;
	ROM[3367] = 4'b0000;
	ROM[3368] = 4'b0000;
	ROM[3369] = 4'b0000;
	ROM[3370] = 4'b0000;
	ROM[3371] = 4'b0000;
	ROM[3372] = 4'b0000;
	ROM[3373] = 4'b0000;
	ROM[3374] = 4'b0000;
	ROM[3375] = 4'b0000;
	ROM[3376] = 4'b0000;
	ROM[3377] = 4'b0000;
	ROM[3378] = 4'b0000;
	ROM[3379] = 4'b0000;
	ROM[3380] = 4'b0000;
	ROM[3381] = 4'b0000;
	ROM[3382] = 4'b0000;
	ROM[3383] = 4'b0000;
	ROM[3384] = 4'b0000;
	ROM[3385] = 4'b0000;
	ROM[3386] = 4'b0000;
	ROM[3387] = 4'b0000;
	ROM[3388] = 4'b0000;
	ROM[3389] = 4'b0000;
	ROM[3390] = 4'b0000;
	ROM[3391] = 4'b0000;
	ROM[3392] = 4'b0000;
	ROM[3393] = 4'b0000;
	ROM[3394] = 4'b0000;
	ROM[3395] = 4'b0000;
	ROM[3396] = 4'b0000;
	ROM[3397] = 4'b0000;
	ROM[3398] = 4'b0000;
	ROM[3399] = 4'b0000;
	ROM[3400] = 4'b0000;
	ROM[3401] = 4'b0000;
	ROM[3402] = 4'b0000;
	ROM[3403] = 4'b0000;
	ROM[3404] = 4'b0000;
	ROM[3405] = 4'b0000;
	ROM[3406] = 4'b0000;
	ROM[3407] = 4'b0000;
	ROM[3408] = 4'b0000;
	ROM[3409] = 4'b0000;
	ROM[3410] = 4'b0000;
	ROM[3411] = 4'b0000;
	ROM[3412] = 4'b0000;
	ROM[3413] = 4'b0000;
	ROM[3414] = 4'b0000;
	ROM[3415] = 4'b0000;
	ROM[3416] = 4'b0000;
	ROM[3417] = 4'b0000;
	ROM[3418] = 4'b0000;
	ROM[3419] = 4'b0000;
	ROM[3420] = 4'b0000;
	ROM[3421] = 4'b0000;
	ROM[3422] = 4'b0000;
	ROM[3423] = 4'b0000;
	ROM[3424] = 4'b0000;
	ROM[3425] = 4'b0000;
	ROM[3426] = 4'b0000;
	ROM[3427] = 4'b0000;
	ROM[3428] = 4'b0000;
	ROM[3429] = 4'b0000;
	ROM[3430] = 4'b0000;
	ROM[3431] = 4'b0000;
	ROM[3432] = 4'b0000;
	ROM[3433] = 4'b0000;
	ROM[3434] = 4'b0000;
	ROM[3435] = 4'b0000;
	ROM[3436] = 4'b0000;
	ROM[3437] = 4'b0000;
	ROM[3438] = 4'b0000;
	ROM[3439] = 4'b0000;
	ROM[3440] = 4'b0000;
	ROM[3441] = 4'b0000;
	ROM[3442] = 4'b0000;
	ROM[3443] = 4'b0000;
	ROM[3444] = 4'b0000;
	ROM[3445] = 4'b0000;
	ROM[3446] = 4'b0000;
	ROM[3447] = 4'b0000;
	ROM[3448] = 4'b0000;
	ROM[3449] = 4'b0000;
	ROM[3450] = 4'b0000;
	ROM[3451] = 4'b0000;
	ROM[3452] = 4'b0000;
	ROM[3453] = 4'b0000;
	ROM[3454] = 4'b0000;
	ROM[3455] = 4'b0000;
	ROM[3456] = 4'b0000;
	ROM[3457] = 4'b0000;
	ROM[3458] = 4'b0000;
	ROM[3459] = 4'b0000;
	ROM[3460] = 4'b0000;
	ROM[3461] = 4'b0000;
	ROM[3462] = 4'b0000;
	ROM[3463] = 4'b0000;
	ROM[3464] = 4'b0000;
	ROM[3465] = 4'b0000;
	ROM[3466] = 4'b0000;
	ROM[3467] = 4'b0000;
	ROM[3468] = 4'b0000;
	ROM[3469] = 4'b0000;
	ROM[3470] = 4'b0000;
	ROM[3471] = 4'b0000;
	ROM[3472] = 4'b0000;
	ROM[3473] = 4'b0000;
	ROM[3474] = 4'b0000;
	ROM[3475] = 4'b0000;
	ROM[3476] = 4'b0000;
	ROM[3477] = 4'b0000;
	ROM[3478] = 4'b0000;
	ROM[3479] = 4'b0000;
	ROM[3480] = 4'b0000;
	ROM[3481] = 4'b0000;
	ROM[3482] = 4'b0000;
	ROM[3483] = 4'b0000;
	ROM[3484] = 4'b0000;
	ROM[3485] = 4'b0000;
	ROM[3486] = 4'b0000;
	ROM[3487] = 4'b0000;
	ROM[3488] = 4'b0000;
	ROM[3489] = 4'b0000;
	ROM[3490] = 4'b0000;
	ROM[3491] = 4'b0000;
	ROM[3492] = 4'b0000;
	ROM[3493] = 4'b0000;
	ROM[3494] = 4'b0000;
	ROM[3495] = 4'b0000;
	ROM[3496] = 4'b0000;
	ROM[3497] = 4'b0000;
	ROM[3498] = 4'b0000;
	ROM[3499] = 4'b0000;
	ROM[3500] = 4'b0000;
	ROM[3501] = 4'b0000;
	ROM[3502] = 4'b0000;
	ROM[3503] = 4'b0000;
	ROM[3504] = 4'b0000;
	ROM[3505] = 4'b0000;
	ROM[3506] = 4'b0000;
	ROM[3507] = 4'b0000;
	ROM[3508] = 4'b0000;
	ROM[3509] = 4'b0000;
	ROM[3510] = 4'b0000;
	ROM[3511] = 4'b0000;
	ROM[3512] = 4'b0000;
	ROM[3513] = 4'b0000;
	ROM[3514] = 4'b0000;
	ROM[3515] = 4'b0000;
	ROM[3516] = 4'b0000;
	ROM[3517] = 4'b0000;
	ROM[3518] = 4'b0000;
	ROM[3519] = 4'b0000;
	ROM[3520] = 4'b0000;
	ROM[3521] = 4'b0000;
	ROM[3522] = 4'b0000;
	ROM[3523] = 4'b0000;
	ROM[3524] = 4'b0000;
	ROM[3525] = 4'b0000;
	ROM[3526] = 4'b0000;
	ROM[3527] = 4'b0000;
	ROM[3528] = 4'b0000;
	ROM[3529] = 4'b0000;
	ROM[3530] = 4'b0000;
	ROM[3531] = 4'b0000;
	ROM[3532] = 4'b0000;
	ROM[3533] = 4'b0000;
	ROM[3534] = 4'b0000;
	ROM[3535] = 4'b0000;
	ROM[3536] = 4'b0000;
	ROM[3537] = 4'b0000;
	ROM[3538] = 4'b0000;
	ROM[3539] = 4'b0000;
	ROM[3540] = 4'b0000;
	ROM[3541] = 4'b0000;
	ROM[3542] = 4'b0000;
	ROM[3543] = 4'b0000;
	ROM[3544] = 4'b0000;
	ROM[3545] = 4'b0000;
	ROM[3546] = 4'b0000;
	ROM[3547] = 4'b0000;
	ROM[3548] = 4'b0000;
	ROM[3549] = 4'b0000;
	ROM[3550] = 4'b0000;
	ROM[3551] = 4'b0000;
	ROM[3552] = 4'b0000;
	ROM[3553] = 4'b0000;
	ROM[3554] = 4'b0000;
	ROM[3555] = 4'b0000;
	ROM[3556] = 4'b0000;
	ROM[3557] = 4'b0000;
	ROM[3558] = 4'b0000;
	ROM[3559] = 4'b0000;
	ROM[3560] = 4'b0000;
	ROM[3561] = 4'b0000;
	ROM[3562] = 4'b0000;
	ROM[3563] = 4'b0000;
	ROM[3564] = 4'b0000;
	ROM[3565] = 4'b0000;
	ROM[3566] = 4'b0000;
	ROM[3567] = 4'b0000;
	ROM[3568] = 4'b0000;
	ROM[3569] = 4'b0000;
	ROM[3570] = 4'b0000;
	ROM[3571] = 4'b0000;
	ROM[3572] = 4'b0000;
	ROM[3573] = 4'b0000;
	ROM[3574] = 4'b0000;
	ROM[3575] = 4'b0000;
	ROM[3576] = 4'b0000;
	ROM[3577] = 4'b0000;
	ROM[3578] = 4'b0000;
	ROM[3579] = 4'b0000;
	ROM[3580] = 4'b0000;
	ROM[3581] = 4'b0000;
	ROM[3582] = 4'b0000;
	ROM[3583] = 4'b0000;
	ROM[3584] = 4'b0000;
	ROM[3585] = 4'b0000;
	ROM[3586] = 4'b0000;
	ROM[3587] = 4'b0000;
	ROM[3588] = 4'b0000;
	ROM[3589] = 4'b0000;
	ROM[3590] = 4'b0000;
	ROM[3591] = 4'b0000;
	ROM[3592] = 4'b0000;
	ROM[3593] = 4'b0000;
	ROM[3594] = 4'b0000;
	ROM[3595] = 4'b0000;
	ROM[3596] = 4'b0000;
	ROM[3597] = 4'b0000;
	ROM[3598] = 4'b0000;
	ROM[3599] = 4'b0000;
	ROM[3600] = 4'b0000;
	ROM[3601] = 4'b0000;
	ROM[3602] = 4'b0000;
	ROM[3603] = 4'b0000;
	ROM[3604] = 4'b0000;
	ROM[3605] = 4'b0000;
	ROM[3606] = 4'b0000;
	ROM[3607] = 4'b0000;
	ROM[3608] = 4'b0000;
	ROM[3609] = 4'b0000;
	ROM[3610] = 4'b0000;
	ROM[3611] = 4'b0000;
	ROM[3612] = 4'b0000;
	ROM[3613] = 4'b0000;
	ROM[3614] = 4'b0000;
	ROM[3615] = 4'b0000;
	ROM[3616] = 4'b0000;
	ROM[3617] = 4'b0000;
	ROM[3618] = 4'b0000;
	ROM[3619] = 4'b0000;
	ROM[3620] = 4'b0000;
	ROM[3621] = 4'b0000;
	ROM[3622] = 4'b0000;
	ROM[3623] = 4'b0000;
	ROM[3624] = 4'b0000;
	ROM[3625] = 4'b0000;
	ROM[3626] = 4'b0000;
	ROM[3627] = 4'b0000;
	ROM[3628] = 4'b0000;
	ROM[3629] = 4'b0000;
	ROM[3630] = 4'b0000;
	ROM[3631] = 4'b0000;
	ROM[3632] = 4'b0000;
	ROM[3633] = 4'b0000;
	ROM[3634] = 4'b0000;
	ROM[3635] = 4'b0000;
	ROM[3636] = 4'b0000;
	ROM[3637] = 4'b0000;
	ROM[3638] = 4'b0000;
	ROM[3639] = 4'b0000;
	ROM[3640] = 4'b0000;
	ROM[3641] = 4'b0000;
	ROM[3642] = 4'b0000;
	ROM[3643] = 4'b0000;
	ROM[3644] = 4'b0000;
	ROM[3645] = 4'b0000;
	ROM[3646] = 4'b0000;
	ROM[3647] = 4'b0000;
	ROM[3648] = 4'b0000;
	ROM[3649] = 4'b0000;
	ROM[3650] = 4'b0000;
	ROM[3651] = 4'b0000;
	ROM[3652] = 4'b0000;
	ROM[3653] = 4'b0000;
	ROM[3654] = 4'b0000;
	ROM[3655] = 4'b0000;
	ROM[3656] = 4'b0000;
	ROM[3657] = 4'b0000;
	ROM[3658] = 4'b0000;
	ROM[3659] = 4'b0000;
	ROM[3660] = 4'b0000;
	ROM[3661] = 4'b0000;
	ROM[3662] = 4'b0000;
	ROM[3663] = 4'b0000;
	ROM[3664] = 4'b0000;
	ROM[3665] = 4'b0000;
	ROM[3666] = 4'b0000;
	ROM[3667] = 4'b0000;
	ROM[3668] = 4'b0000;
	ROM[3669] = 4'b0000;
	ROM[3670] = 4'b0000;
	ROM[3671] = 4'b0000;
	ROM[3672] = 4'b0000;
	ROM[3673] = 4'b0000;
	ROM[3674] = 4'b0000;
	ROM[3675] = 4'b0000;
	ROM[3676] = 4'b0000;
	ROM[3677] = 4'b0000;
	ROM[3678] = 4'b0000;
	ROM[3679] = 4'b0000;
	ROM[3680] = 4'b0000;
	ROM[3681] = 4'b0000;
	ROM[3682] = 4'b0000;
	ROM[3683] = 4'b0000;
	ROM[3684] = 4'b0000;
	ROM[3685] = 4'b0000;
	ROM[3686] = 4'b0000;
	ROM[3687] = 4'b0000;
	ROM[3688] = 4'b0000;
	ROM[3689] = 4'b0000;
	ROM[3690] = 4'b0000;
	ROM[3691] = 4'b0000;
	ROM[3692] = 4'b0000;
	ROM[3693] = 4'b0000;
	ROM[3694] = 4'b0000;
	ROM[3695] = 4'b0000;
	ROM[3696] = 4'b0000;
	ROM[3697] = 4'b0000;
	ROM[3698] = 4'b0000;
	ROM[3699] = 4'b0000;
	ROM[3700] = 4'b0000;
	ROM[3701] = 4'b0000;
	ROM[3702] = 4'b0000;
	ROM[3703] = 4'b0000;
	ROM[3704] = 4'b0000;
	ROM[3705] = 4'b0000;
	ROM[3706] = 4'b0000;
	ROM[3707] = 4'b0000;
	ROM[3708] = 4'b0000;
	ROM[3709] = 4'b0000;
	ROM[3710] = 4'b0000;
	ROM[3711] = 4'b0000;
	ROM[3712] = 4'b0000;
	ROM[3713] = 4'b0000;
	ROM[3714] = 4'b0000;
	ROM[3715] = 4'b0000;
	ROM[3716] = 4'b0000;
	ROM[3717] = 4'b0000;
	ROM[3718] = 4'b0000;
	ROM[3719] = 4'b0000;
	ROM[3720] = 4'b0000;
	ROM[3721] = 4'b0000;
	ROM[3722] = 4'b0000;
	ROM[3723] = 4'b0000;
	ROM[3724] = 4'b0000;
	ROM[3725] = 4'b0000;
	ROM[3726] = 4'b0000;
	ROM[3727] = 4'b0000;
	ROM[3728] = 4'b0000;
	ROM[3729] = 4'b0000;
	ROM[3730] = 4'b0000;
	ROM[3731] = 4'b0000;
	ROM[3732] = 4'b0000;
	ROM[3733] = 4'b0000;
	ROM[3734] = 4'b0000;
	ROM[3735] = 4'b0000;
	ROM[3736] = 4'b0000;
	ROM[3737] = 4'b0000;
	ROM[3738] = 4'b0000;
	ROM[3739] = 4'b0000;
	ROM[3740] = 4'b0000;
	ROM[3741] = 4'b0000;
	ROM[3742] = 4'b0000;
	ROM[3743] = 4'b0000;
	ROM[3744] = 4'b0000;
	ROM[3745] = 4'b0000;
	ROM[3746] = 4'b0000;
	ROM[3747] = 4'b0000;
	ROM[3748] = 4'b0000;
	ROM[3749] = 4'b0000;
	ROM[3750] = 4'b0000;
	ROM[3751] = 4'b0000;
	ROM[3752] = 4'b0000;
	ROM[3753] = 4'b0000;
	ROM[3754] = 4'b0000;
	ROM[3755] = 4'b0000;
	ROM[3756] = 4'b0000;
	ROM[3757] = 4'b0000;
	ROM[3758] = 4'b0000;
	ROM[3759] = 4'b0000;
	ROM[3760] = 4'b0000;
	ROM[3761] = 4'b0000;
	ROM[3762] = 4'b0000;
	ROM[3763] = 4'b0000;
	ROM[3764] = 4'b0000;
	ROM[3765] = 4'b0000;
	ROM[3766] = 4'b0000;
	ROM[3767] = 4'b0000;
	ROM[3768] = 4'b0000;
	ROM[3769] = 4'b0000;
	ROM[3770] = 4'b0000;
	ROM[3771] = 4'b0000;
	ROM[3772] = 4'b0000;
	ROM[3773] = 4'b0000;
	ROM[3774] = 4'b0000;
	ROM[3775] = 4'b0000;
	ROM[3776] = 4'b0000;
	ROM[3777] = 4'b0000;
	ROM[3778] = 4'b0000;
	ROM[3779] = 4'b0000;
	ROM[3780] = 4'b0000;
	ROM[3781] = 4'b0000;
	ROM[3782] = 4'b0000;
	ROM[3783] = 4'b0000;
	ROM[3784] = 4'b0000;
	ROM[3785] = 4'b0000;
	ROM[3786] = 4'b0000;
	ROM[3787] = 4'b0000;
	ROM[3788] = 4'b0000;
	ROM[3789] = 4'b0000;
	ROM[3790] = 4'b0000;
	ROM[3791] = 4'b0000;
	ROM[3792] = 4'b0000;
	ROM[3793] = 4'b0000;
	ROM[3794] = 4'b0000;
	ROM[3795] = 4'b0000;
	ROM[3796] = 4'b0000;
	ROM[3797] = 4'b0000;
	ROM[3798] = 4'b0000;
	ROM[3799] = 4'b0000;
	ROM[3800] = 4'b0000;
	ROM[3801] = 4'b0000;
	ROM[3802] = 4'b0000;
	ROM[3803] = 4'b0000;
	ROM[3804] = 4'b0000;
	ROM[3805] = 4'b0000;
	ROM[3806] = 4'b0000;
	ROM[3807] = 4'b0000;
	ROM[3808] = 4'b0000;
	ROM[3809] = 4'b0000;
	ROM[3810] = 4'b0000;
	ROM[3811] = 4'b0000;
	ROM[3812] = 4'b0000;
	ROM[3813] = 4'b0000;
	ROM[3814] = 4'b0000;
	ROM[3815] = 4'b0000;
	ROM[3816] = 4'b0000;
	ROM[3817] = 4'b0000;
	ROM[3818] = 4'b0000;
	ROM[3819] = 4'b0000;
	ROM[3820] = 4'b0000;
	ROM[3821] = 4'b0000;
	ROM[3822] = 4'b0000;
	ROM[3823] = 4'b0000;
	ROM[3824] = 4'b0000;
	ROM[3825] = 4'b0000;
	ROM[3826] = 4'b0000;
	ROM[3827] = 4'b0000;
	ROM[3828] = 4'b0000;
	ROM[3829] = 4'b0000;
	ROM[3830] = 4'b0000;
	ROM[3831] = 4'b0000;
	ROM[3832] = 4'b0000;
	ROM[3833] = 4'b0000;
	ROM[3834] = 4'b0000;
	ROM[3835] = 4'b0000;
	ROM[3836] = 4'b0000;
	ROM[3837] = 4'b0000;
	ROM[3838] = 4'b0000;
	ROM[3839] = 4'b0000;
	ROM[3840] = 4'b0000;
	ROM[3841] = 4'b0000;
	ROM[3842] = 4'b0000;
	ROM[3843] = 4'b0000;
	ROM[3844] = 4'b0000;
	ROM[3845] = 4'b0000;
	ROM[3846] = 4'b0000;
	ROM[3847] = 4'b0000;
	ROM[3848] = 4'b0000;
	ROM[3849] = 4'b0000;
	ROM[3850] = 4'b0000;
	ROM[3851] = 4'b0000;
	ROM[3852] = 4'b0000;
	ROM[3853] = 4'b0000;
	ROM[3854] = 4'b0000;
	ROM[3855] = 4'b0000;
	ROM[3856] = 4'b0000;
	ROM[3857] = 4'b0000;
	ROM[3858] = 4'b0000;
	ROM[3859] = 4'b0000;
	ROM[3860] = 4'b0000;
	ROM[3861] = 4'b0000;
	ROM[3862] = 4'b0000;
	ROM[3863] = 4'b0000;
	ROM[3864] = 4'b0000;
	ROM[3865] = 4'b0000;
	ROM[3866] = 4'b0000;
	ROM[3867] = 4'b0000;
	ROM[3868] = 4'b0000;
	ROM[3869] = 4'b0000;
	ROM[3870] = 4'b0000;
	ROM[3871] = 4'b0000;
	ROM[3872] = 4'b0000;
	ROM[3873] = 4'b0000;
	ROM[3874] = 4'b0000;
	ROM[3875] = 4'b0000;
	ROM[3876] = 4'b0000;
	ROM[3877] = 4'b0000;
	ROM[3878] = 4'b0000;
	ROM[3879] = 4'b0000;
	ROM[3880] = 4'b0000;
	ROM[3881] = 4'b0000;
	ROM[3882] = 4'b0000;
	ROM[3883] = 4'b0000;
	ROM[3884] = 4'b0000;
	ROM[3885] = 4'b0000;
	ROM[3886] = 4'b0000;
	ROM[3887] = 4'b0000;
	ROM[3888] = 4'b0000;
	ROM[3889] = 4'b0000;
	ROM[3890] = 4'b0000;
	ROM[3891] = 4'b0000;
	ROM[3892] = 4'b0000;
	ROM[3893] = 4'b0000;
	ROM[3894] = 4'b0000;
	ROM[3895] = 4'b0000;
	ROM[3896] = 4'b0000;
	ROM[3897] = 4'b0000;
	ROM[3898] = 4'b0000;
	ROM[3899] = 4'b0000;
	ROM[3900] = 4'b0000;
	ROM[3901] = 4'b0000;
	ROM[3902] = 4'b0000;
	ROM[3903] = 4'b0000;
	ROM[3904] = 4'b0000;
	ROM[3905] = 4'b0000;
	ROM[3906] = 4'b0000;
	ROM[3907] = 4'b0000;
	ROM[3908] = 4'b0000;
	ROM[3909] = 4'b0000;
	ROM[3910] = 4'b0000;
	ROM[3911] = 4'b0000;
	ROM[3912] = 4'b0000;
	ROM[3913] = 4'b0000;
	ROM[3914] = 4'b0000;
	ROM[3915] = 4'b0000;
	ROM[3916] = 4'b0000;
	ROM[3917] = 4'b0000;
	ROM[3918] = 4'b0000;
	ROM[3919] = 4'b0000;
	ROM[3920] = 4'b0000;
	ROM[3921] = 4'b0000;
	ROM[3922] = 4'b0000;
	ROM[3923] = 4'b0000;
	ROM[3924] = 4'b0000;
	ROM[3925] = 4'b0000;
	ROM[3926] = 4'b0000;
	ROM[3927] = 4'b0000;
	ROM[3928] = 4'b0000;
	ROM[3929] = 4'b0000;
	ROM[3930] = 4'b0000;
	ROM[3931] = 4'b0000;
	ROM[3932] = 4'b0000;
	ROM[3933] = 4'b0000;
	ROM[3934] = 4'b0000;
	ROM[3935] = 4'b0000;
	ROM[3936] = 4'b0000;
	ROM[3937] = 4'b0000;
	ROM[3938] = 4'b0000;
	ROM[3939] = 4'b0000;
	ROM[3940] = 4'b0000;
	ROM[3941] = 4'b0000;
	ROM[3942] = 4'b0000;
	ROM[3943] = 4'b0000;
	ROM[3944] = 4'b0000;
	ROM[3945] = 4'b0000;
	ROM[3946] = 4'b0000;
	ROM[3947] = 4'b0000;
	ROM[3948] = 4'b0000;
	ROM[3949] = 4'b0000;
	ROM[3950] = 4'b0000;
	ROM[3951] = 4'b0000;
	ROM[3952] = 4'b0000;
	ROM[3953] = 4'b0000;
	ROM[3954] = 4'b0000;
	ROM[3955] = 4'b0000;
	ROM[3956] = 4'b0000;
	ROM[3957] = 4'b0000;
	ROM[3958] = 4'b0000;
	ROM[3959] = 4'b0000;
	ROM[3960] = 4'b0000;
	ROM[3961] = 4'b0000;
	ROM[3962] = 4'b0000;
	ROM[3963] = 4'b0000;
	ROM[3964] = 4'b0000;
	ROM[3965] = 4'b0000;
	ROM[3966] = 4'b0000;
	ROM[3967] = 4'b0000;
	ROM[3968] = 4'b0000;
	ROM[3969] = 4'b0000;
	ROM[3970] = 4'b0000;
	ROM[3971] = 4'b0000;
	ROM[3972] = 4'b0000;
	ROM[3973] = 4'b0000;
	ROM[3974] = 4'b0000;
	ROM[3975] = 4'b0000;
	ROM[3976] = 4'b0000;
	ROM[3977] = 4'b0000;
	ROM[3978] = 4'b0000;
	ROM[3979] = 4'b0000;
	ROM[3980] = 4'b0000;
	ROM[3981] = 4'b0000;
	ROM[3982] = 4'b0000;
	ROM[3983] = 4'b0000;
	ROM[3984] = 4'b0000;
	ROM[3985] = 4'b0000;
	ROM[3986] = 4'b0000;
	ROM[3987] = 4'b0000;
	ROM[3988] = 4'b0000;
	ROM[3989] = 4'b0000;
	ROM[3990] = 4'b0000;
	ROM[3991] = 4'b0000;
	ROM[3992] = 4'b0000;
	ROM[3993] = 4'b0000;
	ROM[3994] = 4'b0000;
	ROM[3995] = 4'b0000;
	ROM[3996] = 4'b0000;
	ROM[3997] = 4'b0000;
	ROM[3998] = 4'b0000;
	ROM[3999] = 4'b0000;
	ROM[4000] = 4'b0000;
	ROM[4001] = 4'b0000;
	ROM[4002] = 4'b0000;
	ROM[4003] = 4'b0000;
	ROM[4004] = 4'b0000;
	ROM[4005] = 4'b0000;
	ROM[4006] = 4'b0000;
	ROM[4007] = 4'b0000;
	ROM[4008] = 4'b0000;
	ROM[4009] = 4'b0000;
	ROM[4010] = 4'b0000;
	ROM[4011] = 4'b0000;
	ROM[4012] = 4'b0000;
	ROM[4013] = 4'b0000;
	ROM[4014] = 4'b0000;
	ROM[4015] = 4'b0000;
	ROM[4016] = 4'b0000;
	ROM[4017] = 4'b0000;
	ROM[4018] = 4'b0000;
	ROM[4019] = 4'b0000;
	ROM[4020] = 4'b0000;
	ROM[4021] = 4'b0000;
	ROM[4022] = 4'b0000;
	ROM[4023] = 4'b0000;
	ROM[4024] = 4'b0000;
	ROM[4025] = 4'b0000;
	ROM[4026] = 4'b0000;
	ROM[4027] = 4'b0000;
	ROM[4028] = 4'b0000;
	ROM[4029] = 4'b0000;
	ROM[4030] = 4'b0000;
	ROM[4031] = 4'b0000;
	ROM[4032] = 4'b0000;
	ROM[4033] = 4'b0000;
	ROM[4034] = 4'b0000;
	ROM[4035] = 4'b0000;
	ROM[4036] = 4'b0000;
	ROM[4037] = 4'b0000;
	ROM[4038] = 4'b0000;
	ROM[4039] = 4'b0000;
	ROM[4040] = 4'b0000;
	ROM[4041] = 4'b0000;
	ROM[4042] = 4'b0000;
	ROM[4043] = 4'b0000;
	ROM[4044] = 4'b0000;
	ROM[4045] = 4'b0000;
	ROM[4046] = 4'b0000;
	ROM[4047] = 4'b0000;
	ROM[4048] = 4'b0000;
	ROM[4049] = 4'b0000;
	ROM[4050] = 4'b0000;
	ROM[4051] = 4'b0000;
	ROM[4052] = 4'b0000;
	ROM[4053] = 4'b0000;
	ROM[4054] = 4'b0000;
	ROM[4055] = 4'b0000;
	ROM[4056] = 4'b0000;
	ROM[4057] = 4'b0000;
	ROM[4058] = 4'b0000;
	ROM[4059] = 4'b0000;
	ROM[4060] = 4'b0000;
	ROM[4061] = 4'b0000;
	ROM[4062] = 4'b0000;
	ROM[4063] = 4'b0000;
	ROM[4064] = 4'b0000;
	ROM[4065] = 4'b0000;
	ROM[4066] = 4'b0000;
	ROM[4067] = 4'b0000;
	ROM[4068] = 4'b0000;
	ROM[4069] = 4'b0000;
	ROM[4070] = 4'b0000;
	ROM[4071] = 4'b0000;
	ROM[4072] = 4'b0000;
	ROM[4073] = 4'b0000;
	ROM[4074] = 4'b0000;
	ROM[4075] = 4'b0000;
	ROM[4076] = 4'b0000;
	ROM[4077] = 4'b0000;
	ROM[4078] = 4'b0000;
	ROM[4079] = 4'b0000;
	ROM[4080] = 4'b0000;
	ROM[4081] = 4'b0000;
	ROM[4082] = 4'b0000;
	ROM[4083] = 4'b0000;
	ROM[4084] = 4'b0000;
	ROM[4085] = 4'b0000;
	ROM[4086] = 4'b0000;
	ROM[4087] = 4'b0000;
	ROM[4088] = 4'b0000;
	ROM[4089] = 4'b0000;
	ROM[4090] = 4'b0000;
	ROM[4091] = 4'b0000;
	ROM[4092] = 4'b0000;
	ROM[4093] = 4'b0000;
	ROM[4094] = 4'b0000;
	ROM[4095] = 4'b0000;
end

always @(*) begin
    {noteup, notedown} = ROM[addr];
end

endmodule
